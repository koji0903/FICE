//  file name   ... ../../../_library/ice_top_SS3rd_V1.0.35.v
//  top module  ... ../../../_library/ice_top_SS3rd_V1.0.35.v ICE_TOP
//  version     ... V1.0.35
//  designer    ... T.Tsunoda
//  refer to    ... make_chip.para

module ICE_TOP (
  CLK30MHZ_GB ,A19 ,A18 ,A17 ,A16 ,A15 ,A14 ,A13 ,A12 ,A11 ,A10
 ,A9 ,A8 ,A7 ,A6 ,A5 ,A4 ,A3 ,A2 ,DW37 ,DW29
 ,PA13 ,DW36 ,DW28 ,PA12 ,DW35 ,DW27 ,DW19 ,PA11 ,DW34 ,DW26
 ,DW18 ,PA10 ,DW33 ,DW25 ,DW17 ,DDIS ,DW32 ,DW24 ,DW16 ,DW31
 ,DW23 ,DW15 ,DW30 ,DW22 ,DW14 ,DW21 ,DW13 ,ALT1 ,DW20 ,DW12
 ,DW11 ,DW10 ,DW9 ,PA5 ,PC1 ,DW8 ,PA4 ,PC0 ,DW7 ,DIS
 ,PA3 ,DW6 ,PA2 ,DW5 ,DW4 ,DW3 ,DW2 ,DW1 ,MA9 ,DW0
 ,MA8 ,BEU2 ,MA12 ,BEU1 ,MA11 ,BEU0 ,MA10 ,READ ,MRG00 ,MRG01
 ,MRG10 ,MRG11 ,MRG12 ,WWR ,CLKSEL1 ,RDCLKP1 ,FCLK ,PA19 ,PC11 ,PROGI
 ,USBA1 ,CER ,MA2 ,SER ,CE0 ,AF6 ,DA4 ,CE1 ,AF7 ,DA5
 ,EXA ,WED ,EXCH ,MDW0 ,FLMD0 ,SELRO1 ,BRSAM ,ICEWAITMEM ,ICENOECC ,ICEFLERR
 ,RO137 ,RO129 ,EXMA3 ,RO136 ,RO128 ,EXMA2 ,RO135 ,RO127 ,RO119 ,EXMA1
 ,RO134 ,RO126 ,RO118 ,EXMA0 ,RO133 ,RO125 ,RO117 ,RO037 ,RO029 ,RO132
 ,RO124 ,RO116 ,RO036 ,RO028 ,RO131 ,RO123 ,RO115 ,RO035 ,RO027 ,RO019
 ,RO130 ,RO122 ,RO114 ,RO034 ,RO026 ,RO018 ,RO121 ,RO113 ,RO033 ,RO025
 ,RO017 ,RO120 ,RO112 ,RO032 ,RO024 ,RO016 ,RO111 ,RO031 ,RO023 ,RO015
 ,RO110 ,RO030 ,RO022 ,RO014 ,RO19 ,RO18 ,RO17 ,RO09 ,RO16 ,RO08
 ,RO15 ,RO07 ,RO14 ,RO06 ,RO13 ,RO05 ,RO12 ,RO04 ,RO11 ,RO03
 ,MDW9 ,RO10 ,RO02 ,MDW8 ,RO021 ,RO013 ,RO020 ,RO012 ,CPURD ,RO011
 ,RO010 ,RO01 ,MDW7 ,RO00 ,MDW6 ,WAITFL2 ,SLFLASH ,TMEMA14 ,GDRAMWR ,CIBPID31
 ,CIBPID23 ,CIBPID15 ,CIBPID30 ,CIBPID22 ,CIBPID14 ,CIBPID29 ,CIBPID28 ,CIBPID27 ,CIBPID19 ,CIBPID26
 ,CIBPID18 ,CIBPID25 ,CIBPID17 ,CIBPID24 ,CIBPID16 ,CIBPID21 ,CIBPID13 ,CIBPID20 ,CIBPID12 ,CIBPID11
 ,CIBPID10 ,CIBPID9 ,CIBPID8 ,CIBPID7 ,CIBPID6 ,CIBPID5 ,CIBPID4 ,CIBPID3 ,CIBPID2 ,CIBPID1
 ,CIBPID0 ,CPUPID31 ,CPUPID23 ,CPUPID15 ,CPUPID30 ,CPUPID22 ,CPUPID14 ,CPUPID29 ,CPUPID28 ,CPUPID27
 ,CPUPID19 ,CPUPID26 ,CPUPID18 ,CPUPID25 ,CPUPID17 ,CPUPID24 ,CPUPID16 ,CPUPID21 ,CPUPID13 ,CPUPID20
 ,CPUPID12 ,CPUPID11 ,CPUPID10 ,CPUPID9 ,CPUPID8 ,CPUPID7 ,CPUPID6 ,CPUPID5 ,CPUPID4 ,CPUPID3
 ,CPUPID2 ,CPUPID1 ,CPUMASK ,CPUPID0 ,EMEMRAMCLK ,ICEIFA31 ,ICEIFA23 ,ICEIFA15 ,ICEIFA30 ,ICEIFA22
 ,ICEIFA14 ,ICEIFA29 ,ICEIFA28 ,ICEIFA27 ,ICEIFA19 ,ICEIFA26 ,ICEIFA18 ,ICEIFA25 ,ICEIFA17 ,ICEIFA24
 ,ICEIFA16 ,ICEIFA21 ,ICEIFA13 ,ICEDOA29 ,ICEIFA20 ,ICEIFA12 ,ICEDOA28 ,ICEIFA11 ,ICEDOA27 ,ICEDOA19
 ,ICEIFA10 ,ICEDOA26 ,ICEDOA18 ,ICEIFA9 ,ICEIFA8 ,ICEIFA7 ,ICEIFA6 ,ICEIFA5 ,ICEDOA9 ,ICEIFA4
 ,ICEDOA8 ,ICEIFA3 ,ICEDOA7 ,ICEIFA2 ,ICEDOA6 ,ICEIFA1 ,ICEDOA5 ,ICEIFA0 ,ICEDOA4 ,ICEDI31
 ,ICEDI23 ,ICEDI15 ,IDADR11 ,ICEDI30 ,ICEDI22 ,ICEDI14 ,IDADR10 ,ICEDI29 ,IDADR25 ,IDADR17
 ,ICEDI28 ,IDADR24 ,IDADR16 ,ICEDI27 ,ICEDI19 ,IDADR31 ,IDADR23 ,IDADR15 ,ICEDI26 ,ICEDI18
 ,IDADR30 ,IDADR22 ,IDADR14 ,ICEDI25 ,ICEDI17 ,IDADR21 ,IDADR13 ,ICEDI24 ,ICEDI16 ,IDADR20
 ,IDADR12 ,ICEDI21 ,ICEDI13 ,ICEDI20 ,ICEDI12 ,ICEDI11 ,ICEDI10 ,ICEDI9 ,IDADR7 ,ICEDI8
 ,IDADR6 ,ICEDI7 ,IDADR5 ,ICEDI6 ,IDADR4 ,ICEDI5 ,IDADR3 ,ICEDI4 ,IDADR2 ,ICEDI3
 ,IDADR1 ,ICEDI2 ,IDADR0 ,ICEDI1 ,ICEDI0 ,ICEWR ,ICEDOP31 ,ICEDOP23 ,ICEDOP15 ,ICEDOP30
 ,ICEDOP22 ,ICEDOP14 ,ICEDOP29 ,ICEDOP28 ,ICEDOP27 ,ICEDOP19 ,ICEDOP26 ,ICEDOP18 ,ICEDOP25 ,ICEDOP17
 ,ICEDOP24 ,ICEDOP16 ,ICEDOP21 ,ICEDOP13 ,ICEDOP20 ,ICEDOP12 ,ICEDOP11 ,ICEDOP10 ,ICEDOP9 ,ICEDOP8
 ,ICEDOP7 ,ICEDOP6 ,ICEDOP5 ,ICEDOP4 ,ICEDOP3 ,ICEDOP2 ,ICEDOP1 ,ICEDOP0 ,ICEDOA31 ,ICEDOA23
 ,ICEDOA15 ,ICEDOA30 ,ICEDOA22 ,ICEDOA14 ,ICEDOA25 ,ICEDOA17 ,ICEDOA24 ,ICEDOA16 ,ICEDOA21 ,ICEDOA13
 ,ICEDOA20 ,ICEDOA12 ,ICEDOA11 ,ICEDOA10 ,ICEDOA3 ,ICEDOA2 ,ICEDOA1 ,ICEDOA0 ,VDDLEV7 ,VDDLEV6
 ,VDDLEV5 ,VDDLEV4 ,VDDLEV3 ,VDDLEV2 ,VDDLEV1 ,VDDLEV0 ,USBIFWR ,ICECSGREGU ,POCRESB ,TARRESB
 ,CPUPRCLK2 ,CPUTMCLK ,CPUTSCLK ,CPURCLK1SEL ,CLK60MHZ ,CLK60MHZLOCK ,CPUMCLK ,CPUSCLK ,CPURCLK1 ,CPURCLK2
 ,CPURCLK3 ,SOFTBRK ,SVINTACK ,STBRELESV ,SVI ,SVMODI ,SVMODIPERI1 ,SVMODIPERI2 ,SVVCOUT7 ,SVVCOUT6
 ,SVVCOUT5 ,SVVCOUT4 ,SVVCOUT3 ,SVVCOUT2 ,SVVCOUT1 ,SVVCOUT0 ,SVMODOPBRK ,IDADR29 ,IDADR28 ,IDADR27
 ,IDADR19 ,IDADR26 ,IDADR18 ,IDADR9 ,IDADR8 ,PERISVIB ,FLSIZE3 ,FLSIZE2 ,FLSIZE1 ,FLSIZE0
 ,RAMSIZE7 ,RAMSIZE6 ,RAMSIZE5 ,RAMSIZE4 ,RAMSIZE3 ,RAMSIZE2 ,RAMSIZE1 ,RAMSIZE0 ,BFSIZE3 ,BFSIZE2
 ,BFSIZE1 ,BFSIZE0 ,BMSIZE3 ,BMSIZE2 ,BMSIZE1 ,BMSIZE0 ,DFSIZE1 ,DFSIZE0 ,SELRAMMA ,SELDFADMA
 ,PSEUDOON31 ,PSEUDOON23 ,PSEUDOON15 ,PSEUDOON30 ,PSEUDOON22 ,PSEUDOON14 ,PSEUDOON29 ,PSEUDOON28 ,PSEUDOON27 ,PSEUDOON19
 ,PSEUDOON26 ,PSEUDOON18 ,PSEUDOON25 ,PSEUDOON17 ,PSEUDOON24 ,PSEUDOON16 ,PSEUDOON21 ,PSEUDOON13 ,PSEUDOON20 ,PSEUDOON12
 ,PSEUDOON11 ,PSEUDOON10 ,PSEUDOON9 ,PSEUDOON8 ,PSEUDOON7 ,PSEUDOON6 ,PSEUDOON5 ,PSEUDOON4 ,PSEUDOON3 ,PSEUDOON2
 ,PSEUDOON1 ,PSEUDOON0 ,PSEUDOANI09 ,PSEUDOANI17 ,PSEUDOANI08 ,PSEUDOANI16 ,PSEUDOANI07 ,PSEUDOANI15 ,PSEUDOANI06 ,PSEUDOANI14
 ,PSEUDOANI05 ,PSEUDOANI13 ,PSEUDOANI04 ,PSEUDOANI12 ,PSEUDOANI03 ,PSEUDOANI11 ,PSEUDOANI02 ,PSEUDOANI10 ,PSEUDOANI01 ,PSEUDOANI00
 ,PSEUDOANI19 ,PSEUDOANI18 ,ICEMSKDBG ,ICEMSKWAIT ,ICEMSKNMI ,ICEMSKTRAP ,ICEMSKWDT ,ICEMSKLVI ,ICEMSKRETRY ,MDR_RAM15
 ,MDR_RAM14 ,MDR_RAM13 ,MDR_RAM12 ,MDR_RAM11 ,MDR_RAM10 ,MDR_RAM9 ,MDR_RAM8 ,MDR_RAM7 ,MDR_RAM6 ,MDR_RAM5
 ,MDR_RAM4 ,MDR_RAM3 ,MDR_RAM2 ,MDR_RAM1 ,MDR_RAM0 ,CPUWR ,WDOP ,SVMOD ,SVMODF ,STAGEADR1
 ,STAGEADR0 ,PCWAITF ,SKIPEXE ,FCHRAM ,FLREAD ,IMDR10 ,FLREADB3 ,FLREADB2 ,FLREADB1 ,FLREADB0
 ,CPURSOUTB ,BASECK ,PREFIX ,WAITEXM ,OCDWAIT ,BRAMEN ,BFA ,BFAEN ,INTACK ,DMAACK
 ,SLEXM ,IDPOP ,MDW10 ,IMDR2 ,SPINC ,SPDEC ,SPREL ,CPUMISAL ,SLMEM ,FLSPMD
 ,STPST ,HLTST ,MA15 ,MA14 ,MA13 ,MA7 ,MA6 ,MA5 ,MA4 ,MA3
 ,MA1 ,MA0 ,MDW15 ,IMDR7 ,MDW14 ,IMDR6 ,MDW13 ,IMDR5 ,MDW12 ,IMDR4
 ,MDW11 ,IMDR3 ,MDW5 ,MDW4 ,MDW3 ,MDW2 ,MDW1 ,PA18 ,PC10 ,PA17
 ,PA16 ,PA15 ,PA14 ,PA9 ,PC5 ,PA8 ,PC4 ,PA7 ,PC3 ,PA6
 ,PC2 ,PC19 ,PC18 ,PC17 ,PC16 ,PC15 ,PC14 ,PC13 ,PC12 ,PC9
 ,PC8 ,PC7 ,PC6 ,IMDR15 ,IMDR14 ,IMDR13 ,IMDR12 ,IMDR11 ,IMDR9 ,IMDR8
 ,IMDR1 ,IMDR0 ,SLBMEM ,SYSRSOUTB ,PONRESB ,CPUPRCLK3 ,LOCKFAIL5 ,LOCKFAIL6 ,LOCKFAIL7 ,LOCKFAIL8
 ,LOCKFAIL9 ,LOCKFAIL10 ,LOCKFAIL11 ,LOCKFAIL12 ,LOCKFAIL20 ,LOCKFAIL13 ,LOCKFAIL21 ,LOCKFAIL14 ,LOCKFAIL22 ,LOCKFAIL30
 ,LOCKFAIL15 ,LOCKFAIL23 ,LOCKFAIL16 ,LOCKFAIL24 ,LOCKFAIL17 ,LOCKFAIL25 ,LOCKFAIL18 ,LOCKFAIL26 ,LOCKFAIL19 ,LOCKFAIL27
 ,LOCKFAIL28 ,LOCKFAIL29 ,IDVER31 ,IDVER23 ,IDVER15 ,IDVER30 ,IDVER22 ,IDVER14 ,IDVER29 ,IDVER28
 ,IDVER27 ,IDVER19 ,IDVER26 ,IDVER18 ,IDVER25 ,IDVER17 ,IDVER24 ,IDVER16 ,IDVER21 ,IDVER13
 ,IDVER20 ,IDVER12 ,IDVER11 ,IDVER10 ,IDVER9 ,IDVER8 ,IDVER7 ,IDVER6 ,IDVER5 ,IDVER4
 ,IDVER3 ,IDVER2 ,IDVER1 ,IDVER0 ,ADDRTD144 ,ADDRTD136 ,ADDRTD128 ,ADDRTD143 ,ADDRTD135 ,ADDRTD127
 ,ADDRTD119 ,ADDRTD142 ,ADDRTD134 ,ADDRTD126 ,ADDRTD118 ,ADDRTD141 ,ADDRTD133 ,ADDRTD125 ,ADDRTD117 ,ADDRTD109
 ,ADDRTD140 ,ADDRTD132 ,ADDRTD124 ,ADDRTD116 ,ADDRTD108 ,ADDRTD139 ,ADDRTD138 ,ADDRTD137 ,ADDRTD129 ,ADDRTD131
 ,ADDRTD123 ,ADDRTD115 ,ADDRTD107 ,ADDRTD130 ,ADDRTD122 ,ADDRTD114 ,ADDRTD106 ,ADDRTD121 ,ADDRTD113 ,ADDRTD105
 ,ADDRTD120 ,ADDRTD112 ,ADDRTD104 ,ADDRTD111 ,ADDRTD103 ,ADDRTD110 ,ADDRTD102 ,ADDRTD101 ,ADDRTD100 ,ADDRTD99
 ,ADDRTD98 ,ADDRTD97 ,ADDRTD89 ,ADDRTD96 ,ADDRTD88 ,ADDRTD95 ,ADDRTD87 ,ADDRTD79 ,ADDRTD94 ,ADDRTD86
 ,ADDRTD78 ,ADDRTD93 ,ADDRTD85 ,ADDRTD77 ,ADDRTD69 ,ADDRTD92 ,ADDRTD84 ,ADDRTD76 ,ADDRTD68 ,ADDRTD91
 ,ADDRTD83 ,ADDRTD75 ,ADDRTD67 ,ADDRTD59 ,ADDRTD90 ,ADDRTD82 ,ADDRTD74 ,ADDRTD66 ,ADDRTD58 ,ADDRTD81
 ,ADDRTD73 ,ADDRTD65 ,ADDRTD57 ,ADDRTD49 ,ADDRTD80 ,ADDRTD72 ,ADDRTD64 ,ADDRTD56 ,ADDRTD48 ,ADDRTD71
 ,ADDRTD63 ,ADDRTD55 ,ADDRTD47 ,ADDRTD39 ,ADDRTD70 ,ADDRTD62 ,ADDRTD54 ,ADDRTD46 ,ADDRTD38 ,ADDRTD61
 ,ADDRTD53 ,ADDRTD45 ,ADDRTD37 ,ADDRTD29 ,ADDRTD60 ,ADDRTD52 ,ADDRTD44 ,ADDRTD36 ,ADDRTD28 ,ADDRTD51
 ,ADDRTD43 ,ADDRTD35 ,ADDRTD27 ,ADDRTD19 ,ADDRTD50 ,ADDRTD42 ,ADDRTD34 ,ADDRTD26 ,ADDRTD18 ,ADDRTD41
 ,ADDRTD33 ,ADDRTD25 ,ADDRTD17 ,ADDRTD40 ,ADDRTD32 ,ADDRTD24 ,ADDRTD16 ,ADDRTD31 ,ADDRTD23 ,ADDRTD15
 ,ADDRTD30 ,ADDRTD22 ,ADDRTD14 ,ADDRTD21 ,ADDRTD13 ,ADDRTD20 ,ADDRTD12 ,ADDRTD11 ,ADDRTD10 ,ADDRTD9
 ,ADDRTD8 ,ADDRTD7 ,ADDRTD6 ,ADDRTD5 ,ADDRTD4 ,ADDRTD3 ,ADDRTD2 ,ADDRTD1 ,ADDRPINRD ,ADDRPINMD
 ,ADDRPINLV ,TP144D3 ,TP136D3 ,TP128D3 ,TP144D2 ,TP136D2 ,TP128D2 ,TP144D1 ,TP136D1 ,TP128D1
 ,TP144D0 ,TP136D0 ,TP128D0 ,TP143D3 ,TP135D3 ,TP127D3 ,TP119D3 ,TP143D2 ,TP135D2 ,TP127D2
 ,TP119D2 ,TP143D1 ,TP135D1 ,TP127D1 ,TP119D1 ,TP143D0 ,TP135D0 ,TP127D0 ,TP119D0 ,TP142D3
 ,TP134D3 ,TP126D3 ,TP118D3 ,TP142D2 ,TP134D2 ,TP126D2 ,TP118D2 ,TP142D1 ,TP134D1 ,TP126D1
 ,TP118D1 ,TP142D0 ,TP134D0 ,TP126D0 ,TP118D0 ,TP141D3 ,TP133D3 ,TP125D3 ,TP117D3 ,TP109D3
 ,TP141D2 ,TP133D2 ,TP125D2 ,TP117D2 ,TP109D2 ,TP141D1 ,TP133D1 ,TP125D1 ,TP117D1 ,TP109D1
 ,TP141D0 ,TP133D0 ,TP125D0 ,TP117D0 ,TP109D0 ,TP140D3 ,TP132D3 ,TP124D3 ,TP116D3 ,TP108D3
 ,TP140D2 ,TP132D2 ,TP124D2 ,TP116D2 ,TP108D2 ,TP140D1 ,TP132D1 ,TP124D1 ,TP116D1 ,TP108D1
 ,TP140D0 ,TP132D0 ,TP124D0 ,TP116D0 ,TP108D0 ,TP139D3 ,TP139D2 ,TP139D1 ,TP139D0 ,TP138D3
 ,TP138D2 ,TP138D1 ,TP138D0 ,TP137D3 ,TP129D3 ,TP137D2 ,TP129D2 ,TP137D1 ,TP129D1 ,TP137D0
 ,TP129D0 ,TP131D3 ,TP123D3 ,TP115D3 ,TP107D3 ,TP131D2 ,TP123D2 ,TP115D2 ,TP107D2 ,TP131D1
 ,TP123D1 ,TP115D1 ,TP107D1 ,TP131D0 ,TP123D0 ,TP115D0 ,TP107D0 ,TP130D3 ,TP122D3 ,TP114D3
 ,TP106D3 ,TP130D2 ,TP122D2 ,TP114D2 ,TP106D2 ,TP130D1 ,TP122D1 ,TP114D1 ,TP106D1 ,TP130D0
 ,TP122D0 ,TP114D0 ,TP106D0 ,TP121D3 ,TP113D3 ,TP105D3 ,TP121D2 ,TP113D2 ,TP105D2 ,TP121D1
 ,TP113D1 ,TP105D1 ,TP121D0 ,TP113D0 ,TP105D0 ,TP120D3 ,TP112D3 ,TP104D3 ,TP120D2 ,TP112D2
 ,TP104D2 ,EROMWRB ,TP120D1 ,TP112D1 ,TP104D1 ,TP120D0 ,TP112D0 ,TP104D0 ,TP111D3 ,TP103D3
 ,TP111D2 ,TP103D2 ,TP111D1 ,TP103D1 ,TP111D0 ,TP103D0 ,TP110D3 ,TP102D3 ,TP110D2 ,TP102D2
 ,TP110D1 ,TP102D1 ,TP110D0 ,TP102D0 ,TP101D3 ,TP101D2 ,TP101D1 ,TP101D0 ,TP100D3 ,TP100D2
 ,TP100D1 ,TP100D0 ,TP99D3 ,TP99D2 ,TP99D1 ,TP99D0 ,TP98D3 ,TP98D2 ,TP98D1 ,TP98D0
 ,TP97D3 ,TP89D3 ,TP97D2 ,TP89D2 ,TP97D1 ,TP89D1 ,TP97D0 ,TP89D0 ,TP96D3 ,TP88D3
 ,TP96D2 ,TP88D2 ,TP96D1 ,TP88D1 ,TP96D0 ,TP88D0 ,TP95D3 ,TP87D3 ,TP79D3 ,TP95D2
 ,TP87D2 ,TP79D2 ,TP95D1 ,TP87D1 ,TP79D1 ,TP95D0 ,TP87D0 ,TP79D0 ,TP94D3 ,TP86D3
 ,TP78D3 ,TP94D2 ,TP86D2 ,TP78D2 ,TP94D1 ,TP86D1 ,TP78D1 ,TP94D0 ,TP86D0 ,TP78D0
 ,TP93D3 ,TP85D3 ,TP77D3 ,TP69D3 ,TP93D2 ,TP85D2 ,TP77D2 ,TP69D2 ,TP93D1 ,TP85D1
 ,TP77D1 ,TP69D1 ,TP93D0 ,TP85D0 ,TP77D0 ,TP69D0 ,TP92D3 ,TP84D3 ,TP76D3 ,TP68D3
 ,TP92D2 ,TP84D2 ,TP76D2 ,TP68D2 ,TP92D1 ,TP84D1 ,TP76D1 ,TP68D1 ,TP92D0 ,TP84D0
 ,TP76D0 ,TP68D0 ,TP91D3 ,TP83D3 ,TP75D3 ,TP67D3 ,TP59D3 ,TP91D2 ,TP83D2 ,TP75D2
 ,TP67D2 ,TP59D2 ,TP91D1 ,TP83D1 ,TP75D1 ,TP67D1 ,TP59D1 ,TP91D0 ,TP83D0 ,TP75D0
 ,TP67D0 ,TP59D0 ,TP90D3 ,TP82D3 ,TP74D3 ,TP66D3 ,TP58D3 ,TP90D2 ,TP82D2 ,TP74D2
 ,TP66D2 ,TP58D2 ,TP90D1 ,TP82D1 ,TP74D1 ,TP66D1 ,TP58D1 ,TP90D0 ,TP82D0 ,TP74D0
 ,TP66D0 ,TP58D0 ,TP81D3 ,TP73D3 ,TP65D3 ,TP57D3 ,TP49D3 ,TP81D2 ,TP73D2 ,TP65D2
 ,TP57D2 ,TP49D2 ,TP81D1 ,TP73D1 ,TP65D1 ,TP57D1 ,TP49D1 ,TP81D0 ,TP73D0 ,TP65D0
 ,TP57D0 ,TP49D0 ,TP80D3 ,TP72D3 ,TP64D3 ,TP56D3 ,TP48D3 ,TP80D2 ,TP72D2 ,TP64D2
 ,TP56D2 ,TP48D2 ,TP80D1 ,TP72D1 ,TP64D1 ,TP56D1 ,TP48D1 ,TP80D0 ,TP72D0 ,TP64D0
 ,TP56D0 ,TP48D0 ,TP71D3 ,TP63D3 ,TP55D3 ,TP47D3 ,TP39D3 ,TP71D2 ,TP63D2 ,TP55D2
 ,TP47D2 ,TP39D2 ,TP71D1 ,TP63D1 ,TP55D1 ,TP47D1 ,TP39D1 ,TP71D0 ,TP63D0 ,TP55D0
 ,TP47D0 ,TP39D0 ,TP70D3 ,TP62D3 ,TP54D3 ,TP46D3 ,TP38D3 ,TP70D2 ,TP62D2 ,TP54D2
 ,TP46D2 ,TP38D2 ,TP70D1 ,TP62D1 ,TP54D1 ,TP46D1 ,TP38D1 ,TP70D0 ,TP62D0 ,TP54D0
 ,TP46D0 ,TP38D0 ,TP61D3 ,TP53D3 ,TP45D3 ,TP37D3 ,TP29D3 ,TP61D2 ,TP53D2 ,TP45D2
 ,TP37D2 ,TP29D2 ,TP61D1 ,TP53D1 ,TP45D1 ,TP37D1 ,TP29D1 ,TP61D0 ,TP53D0 ,TP45D0
 ,TP37D0 ,TP29D0 ,TP60D3 ,TP52D3 ,TP44D3 ,TP36D3 ,TP28D3 ,TP60D2 ,TP52D2 ,TP44D2
 ,TP36D2 ,TP28D2 ,TP60D1 ,TP52D1 ,TP44D1 ,TP36D1 ,TP28D1 ,TP60D0 ,TP52D0 ,TP44D0
 ,TP36D0 ,TP28D0 ,TP51D3 ,TP43D3 ,TP35D3 ,TP27D3 ,TP19D3 ,TP51D2 ,TP43D2 ,TP35D2
 ,TP27D2 ,TP19D2 ,TP51D1 ,TP43D1 ,TP35D1 ,TP27D1 ,TP19D1 ,TP51D0 ,TP43D0 ,TP35D0
 ,TP27D0 ,TP19D0 ,TP50D3 ,TP42D3 ,TP34D3 ,TP26D3 ,TP18D3 ,TP50D2 ,TP42D2 ,TP34D2
 ,TP26D2 ,TP18D2 ,TP50D1 ,TP42D1 ,TP34D1 ,TP26D1 ,TP18D1 ,TP50D0 ,TP42D0 ,TP34D0
 ,TP26D0 ,TP18D0 ,TP41D3 ,TP33D3 ,TP25D3 ,TP17D3 ,TP41D2 ,TP33D2 ,TP25D2 ,TP17D2
 ,TP41D1 ,TP33D1 ,TP25D1 ,TP17D1 ,TP41D0 ,TP33D0 ,TP25D0 ,TP17D0 ,TP40D3 ,TP32D3
 ,TP24D3 ,TP16D3 ,TP40D2 ,TP32D2 ,TP24D2 ,TP16D2 ,TP40D1 ,TP32D1 ,TP24D1 ,TP16D1
 ,TP40D0 ,TP32D0 ,TP24D0 ,TP16D0 ,TP31D3 ,TP23D3 ,TP15D3 ,TP31D2 ,TP23D2 ,TP15D2
 ,TP31D1 ,TP23D1 ,TP15D1 ,TP31D0 ,TP23D0 ,TP15D0 ,TP30D3 ,TP22D3 ,TP14D3 ,TP30D2
 ,TP22D2 ,TP14D2 ,TP30D1 ,TP22D1 ,TP14D1 ,TP30D0 ,TP22D0 ,TP14D0 ,TP21D3 ,TP13D3
 ,TP21D2 ,TP13D2 ,TP21D1 ,TP13D1 ,TP21D0 ,TP13D0 ,TP20D3 ,TP12D3 ,TP20D2 ,TP12D2
 ,TP20D1 ,TP12D1 ,TP20D0 ,TP12D0 ,TP11D3 ,TP11D2 ,TP11D1 ,TP11D0 ,TP10D3 ,TP10D2
 ,TP10D1 ,TP10D0 ,TP9D3 ,TP9D2 ,TP9D1 ,TP9D0 ,TP8D3 ,TP8D2 ,TP8D1 ,TP8D0
 ,TP7D3 ,TP7D2 ,TP7D1 ,TP7D0 ,TP6D3 ,TP6D2 ,TP6D1 ,TP6D0 ,TP5D3 ,TP5D2
 ,TP5D1 ,TP5D0 ,TP4D3 ,TP4D2 ,TP4D1 ,TP4D0 ,TP3D3 ,TP3D2 ,TP3D1 ,TP3D0
 ,TP2D3 ,TP2D2 ,TP2D1 ,TP2D0 ,TP1D3 ,TP1D2 ,TP1D1 ,TP1D0 ,CLK30MHZ ,EROMRDB
 ,EROMCSB ,EROMPA2 ,EROMCLK ,EROMPA17 ,EROMPA16 ,EROMPA15 ,EROMPA14 ,EROMPA13 ,EROMPA12 ,EROMPA11
 ,EROMPA10 ,EROMPA9 ,EROMPD3 ,EROMPA8 ,EROMPD2 ,EROMPA7 ,EROMPD1 ,EROMPA6 ,EROMPD0 ,EROMPA5
 ,EROMPA4 ,EROMPA3 ,EROMPA1 ,EROMPA0 ,RDCLKP1_OUT ,EXA_OUT ,WWR_OUT ,CER_OUT ,SER_OUT ,EXER_OUT
 ,MRG00_OUT ,MRG01_OUT ,MRG10_OUT ,MRG11_OUT ,MRG12_OUT ,DIS_OUT ,READ_OUT ,FCLK_OUT ,PROGI_OUT ,BFA_OUT
 ,EROMPD31 ,EROMPD23 ,EROMPD15 ,EROMPD30 ,EROMPD22 ,EROMPD14 ,EROMPD29 ,EROMPD28 ,EROMPD27 ,EROMPD19
 ,EROMPD26 ,EROMPD18 ,EROMPD25 ,EROMPD17 ,EROMPD24 ,EROMPD16 ,EROMPD21 ,EROMPD13 ,EROMPD20 ,EROMPD12
 ,EROMPD11 ,EROMPD10 ,EROMPD9 ,EROMPD8 ,EROMPD7 ,EROMPD6 ,EROMPD5 ,EROMPD4 ,BTFLG ,TMSPMD
 ,TMBTSEL ,ICETMSPMD ,ICETMBTSEL ,RESB ,USBCLK ,USBRD_B ,USBWR0_B ,USBA21 ,USBA20 ,USBA19
 ,USBA4 ,USBA3 ,USBA2 ,USBWAIT_B ,USBD15 ,USBD14 ,USBD13 ,USBD12 ,USBD11 ,USBD10
 ,USBD9 ,USBD8 ,USBD7 ,USBD6 ,USBD5 ,USBD4 ,USBD3 ,USBD2 ,USBD1 ,USBD0
 ,ICESYSRES_B ,ICECPURES_B ,RESET_B ,EVAOSCMCLK ,EVAOSCRCLK1 ,EVAOSCRCLK2 ,EVAOSCRCLK3 ,TMEMA16 ,TMEMA15 ,TMEMA13
 ,TMEMA12 ,TMEMA11 ,TMEMA10 ,TMEMA9 ,TMEMD3 ,TMEMA8 ,TMEMD2 ,TMEMA7 ,TMEMD1 ,TMEMA6
 ,TMEMD0 ,TMEMA5 ,TMEMA4 ,TMEMA3 ,TMEMA2 ,TMEMA1 ,TMEMA0 ,TMEMCS_B ,TMEMRD_B ,TMEMWR_B
 ,TMEMCLK2 ,TMEMCLK1 ,TMEMCLK0 ,TMEMD107 ,TMEMD106 ,TMEMD105 ,TMEMD104 ,TMEMD103 ,TMEMD102 ,TMEMD101
 ,TMEMD100 ,TMEMD99 ,TMEMD98 ,TMEMD97 ,TMEMD89 ,TMEMD96 ,TMEMD88 ,TMEMD95 ,TMEMD87 ,TMEMD79
 ,TMEMD94 ,TMEMD86 ,TMEMD78 ,TMEMD93 ,TMEMD85 ,TMEMD77 ,TMEMD69 ,TMEMD92 ,TMEMD84 ,TMEMD76
 ,TMEMD68 ,TMEMD91 ,TMEMD83 ,TMEMD75 ,TMEMD67 ,TMEMD59 ,TMEMD90 ,TMEMD82 ,TMEMD74 ,TMEMD66
 ,TMEMD58 ,TMEMD81 ,TMEMD73 ,TMEMD65 ,TMEMD57 ,TMEMD49 ,TMEMD80 ,TMEMD72 ,TMEMD64 ,TMEMD56
 ,TMEMD48 ,TMEMD71 ,TMEMD63 ,TMEMD55 ,TMEMD47 ,TMEMD39 ,TMEMD70 ,TMEMD62 ,TMEMD54 ,TMEMD46
 ,TMEMD38 ,TMEMD61 ,TMEMD53 ,TMEMD45 ,TMEMD37 ,TMEMD29 ,TMEMD60 ,TMEMD52 ,TMEMD44 ,TMEMD36
 ,TMEMD28 ,TMEMD51 ,TMEMD43 ,TMEMD35 ,TMEMD27 ,TMEMD19 ,TMEMD50 ,TMEMD42 ,TMEMD34 ,TMEMD26
 ,TMEMD18 ,TMEMD41 ,TMEMD33 ,TMEMD25 ,TMEMD17 ,TMEMD40 ,TMEMD32 ,TMEMD24 ,TMEMD16 ,TMEMD31
 ,TMEMD23 ,TMEMD15 ,TMEMD30 ,TMEMD22 ,TMEMD14 ,TMEMD21 ,TMEMD13 ,TMEMD20 ,TMEMD12 ,TMEMD11
 ,TMEMD10 ,TMEMD9 ,TMEMD8 ,TMEMD7 ,TMEMD6 ,TMEMD5 ,TMEMD4 ,TCCONNECT_B ,EACONNECT_B ,TVDDON
 ,TVDDSEL ,LEDTVDD_B ,LEDCLOCK_B ,LEDRUN_B ,LEDRESET_B ,LEDSTANDBY_B ,LEDWAIT_B ,DCE0 ,DCLKSEL1 ,DCER
 ,DSER ,DWWR ,DWED ,DMRG00 ,DMRG01 ,DMRG10 ,DMRG11 ,DMRG12 ,DREAD ,AF19
 ,AF18 ,AF17 ,DA13 ,AF16 ,DA12 ,AF15 ,DA11 ,AF14 ,DA10 ,AF13
 ,AF12 ,AF11 ,AF10 ,AF9 ,DA7 ,AF8 ,DA6 ,AF5 ,DA3 ,AF4
 ,DA2 ,AF3 ,DA1 ,AF2 ,DA0 ,AF1 ,AF0 ,DRDCLK ,DRDCLKC1 ,DA9
 ,DA8 ,DRO11 ,DRO10 ,DRO9 ,DRO8 ,DRO7 ,DRO6 ,DRO5 ,DRO4 ,DRO3
 ,DRO2 ,DRO1 ,DRO0 ,DDIS_OUT ,DRDCLKP1_OUT ,DWWR_OUT ,DCER_OUT ,DSER_OUT ,DMRG00_OUT ,DMRG01_OUT
 ,DMRG10_OUT ,DMRG11_OUT ,DMRG12_OUT ,DREAD_OUT ,DFCLK_OUT ,SLDFLASH ,LOCK240FAIL ,CLK240M ,CLK120M
);

  input A19 ,A18 ,A17 ,A16 ,A15 ,A14 ,A13 ,A12 ,A11 ;
  input A10 ,A9 ,A8 ,A7 ,A6 ,A5 ,A4 ,A3 ,A2 ;
  input DW37 ,DW29 ,PA13 ,DW36 ,DW28 ,PA12 ,DW35 ,DW27 ,DW19 ;
  input PA11 ,DW34 ,DW26 ,DW18 ,PA10 ,DW33 ,DW25 ,DW17 ,DDIS ;
  input DW32 ,DW24 ,DW16 ,DW31 ,DW23 ,DW15 ,DW30 ,DW22 ,DW14 ;
  input DW21 ,DW13 ,ALT1 ,DW20 ,DW12 ,DW11 ,DW10 ,DW9 ,PA5 ;
  input PC1 ,DW8 ,PA4 ,PC0 ,DW7 ,DIS ,PA3 ,DW6 ,PA2 ;
  input DW5 ,DW4 ,DW3 ,DW2 ,DW1 ,MA9 ,DW0 ,MA8 ,BEU2 ;
  input MA12 ,BEU1 ,MA11 ,BEU0 ,MA10 ,READ ,MRG00 ,MRG01 ,MRG10 ;
  input MRG11 ,MRG12 ,WWR ,CLKSEL1 ,RDCLKP1 ,FCLK ,PA19 ,PC11 ,PROGI ;
  input USBA1 ,CER ,MA2 ,SER ,CE0 ,AF6 ,DA4 ,CE1 ,AF7 ;
  input DA5 ,EXA ,WED ,EXCH ,MDW0 ,FLMD0 ,SELRO1 ,BRSAM ,EXMA3 ;
  input EXMA2 ,EXMA1 ,EXMA0 ,MDW9 ,MDW8 ,CPURD ,MDW7 ,MDW6 ,SLFLASH ;
  input GDRAMWR ,CIBPID31 ,CIBPID23 ,CIBPID15 ,CIBPID30 ,CIBPID22 ,CIBPID14 ,CIBPID29 ,CIBPID28 ;
  input CIBPID27 ,CIBPID19 ,CIBPID26 ,CIBPID18 ,CIBPID25 ,CIBPID17 ,CIBPID24 ,CIBPID16 ,CIBPID21 ;
  input CIBPID13 ,CIBPID20 ,CIBPID12 ,CIBPID11 ,CIBPID10 ,CIBPID9 ,CIBPID8 ,CIBPID7 ,CIBPID6 ;
  input CIBPID5 ,CIBPID4 ,CIBPID3 ,CIBPID2 ,CIBPID1 ,CIBPID0 ,CPUMASK ,EMEMRAMCLK ,ICEDOA29 ;
  input ICEDOA28 ,ICEDOA27 ,ICEDOA19 ,ICEDOA26 ,ICEDOA18 ,ICEDOA9 ,ICEDOA8 ,ICEDOA7 ,ICEDOA6 ;
  input ICEDOA5 ,ICEDOA4 ,IDADR11 ,IDADR10 ,IDADR25 ,IDADR17 ,IDADR24 ,IDADR16 ,IDADR31 ;
  input IDADR23 ,IDADR15 ,IDADR30 ,IDADR22 ,IDADR14 ,IDADR21 ,IDADR13 ,IDADR20 ,IDADR12 ;
  input IDADR7 ,IDADR6 ,IDADR5 ,IDADR4 ,IDADR3 ,IDADR2 ,IDADR1 ,IDADR0 ,ICEDOP31 ;
  input ICEDOP23 ,ICEDOP15 ,ICEDOP30 ,ICEDOP22 ,ICEDOP14 ,ICEDOP29 ,ICEDOP28 ,ICEDOP27 ,ICEDOP19 ;
  input ICEDOP26 ,ICEDOP18 ,ICEDOP25 ,ICEDOP17 ,ICEDOP24 ,ICEDOP16 ,ICEDOP21 ,ICEDOP13 ,ICEDOP20 ;
  input ICEDOP12 ,ICEDOP11 ,ICEDOP10 ,ICEDOP9 ,ICEDOP8 ,ICEDOP7 ,ICEDOP6 ,ICEDOP5 ,ICEDOP4 ;
  input ICEDOP3 ,ICEDOP2 ,ICEDOP1 ,ICEDOP0 ,ICEDOA31 ,ICEDOA23 ,ICEDOA15 ,ICEDOA30 ,ICEDOA22 ;
  input ICEDOA14 ,ICEDOA25 ,ICEDOA17 ,ICEDOA24 ,ICEDOA16 ,ICEDOA21 ,ICEDOA13 ,ICEDOA20 ,ICEDOA12 ;
  input ICEDOA11 ,ICEDOA10 ,ICEDOA3 ,ICEDOA2 ,ICEDOA1 ,ICEDOA0 ,CPUPRCLK2 ,CPUTMCLK ,CPUTSCLK ;
  input CPURCLK1SEL ,SOFTBRK ,SVINTACK ,IDADR29 ,IDADR28 ,IDADR27 ,IDADR19 ,IDADR26 ,IDADR18 ;
  input IDADR9 ,IDADR8 ,PERISVIB ,CPUWR ,WDOP ,SVMOD ,SVMODF ,STAGEADR1 ,STAGEADR0 ;
  input PCWAITF ,SKIPEXE ,FCHRAM ,FLREAD ,IMDR10 ,FLREADB3 ,FLREADB2 ,FLREADB1 ,FLREADB0 ;
  input CPURSOUTB ,BASECK ,PREFIX ,WAITEXM ,OCDWAIT ,BRAMEN ,BFA ,BFAEN ,INTACK ;
  input DMAACK ,SLEXM ,IDPOP ,MDW10 ,IMDR2 ,SPINC ,SPDEC ,SPREL ,CPUMISAL ;
  input SLMEM ,FLSPMD ,STPST ,HLTST ,MA15 ,MA14 ,MA13 ,MA7 ,MA6 ;
  input MA5 ,MA4 ,MA3 ,MA1 ,MA0 ,MDW15 ,IMDR7 ,MDW14 ,IMDR6 ;
  input MDW13 ,IMDR5 ,MDW12 ,IMDR4 ,MDW11 ,IMDR3 ,MDW5 ,MDW4 ,MDW3 ;
  input MDW2 ,MDW1 ,PA18 ,PC10 ,PA17 ,PA16 ,PA15 ,PA14 ,PA9 ;
  input PC5 ,PA8 ,PC4 ,PA7 ,PC3 ,PA6 ,PC2 ,PC19 ,PC18 ;
  input PC17 ,PC16 ,PC15 ,PC14 ,PC13 ,PC12 ,PC9 ,PC8 ,PC7 ;
  input PC6 ,IMDR15 ,IMDR14 ,IMDR13 ,IMDR12 ,IMDR11 ,IMDR9 ,IMDR8 ,IMDR1 ;
  input IMDR0 ,SLBMEM ,CPUPRCLK3 ,LOCKFAIL5 ,LOCKFAIL6 ,LOCKFAIL7 ,LOCKFAIL8 ,LOCKFAIL9 ,LOCKFAIL10 ;
  input LOCKFAIL11 ,LOCKFAIL12 ,LOCKFAIL20 ,LOCKFAIL13 ,LOCKFAIL21 ,LOCKFAIL14 ,LOCKFAIL22 ,LOCKFAIL30 ,LOCKFAIL15 ;
  input LOCKFAIL23 ,LOCKFAIL16 ,LOCKFAIL24 ,LOCKFAIL17 ,LOCKFAIL25 ,LOCKFAIL18 ,LOCKFAIL26 ,LOCKFAIL19 ,LOCKFAIL27 ;
  input LOCKFAIL28 ,LOCKFAIL29 ,IDVER31 ,IDVER23 ,IDVER15 ,IDVER30 ,IDVER22 ,IDVER14 ,IDVER29 ;
  input IDVER28 ,IDVER27 ,IDVER19 ,IDVER26 ,IDVER18 ,IDVER25 ,IDVER17 ,IDVER24 ,IDVER16 ;
  input IDVER21 ,IDVER13 ,IDVER20 ,IDVER12 ,IDVER11 ,IDVER10 ,IDVER9 ,IDVER8 ,IDVER7 ;
  input IDVER6 ,IDVER5 ,IDVER4 ,IDVER3 ,IDVER2 ,IDVER1 ,IDVER0 ,TP144D3 ,TP136D3 ;
  input TP128D3 ,TP144D2 ,TP136D2 ,TP128D2 ,TP144D1 ,TP136D1 ,TP128D1 ,TP144D0 ,TP136D0 ;
  input TP128D0 ,TP143D3 ,TP135D3 ,TP127D3 ,TP119D3 ,TP143D2 ,TP135D2 ,TP127D2 ,TP119D2 ;
  input TP143D1 ,TP135D1 ,TP127D1 ,TP119D1 ,TP143D0 ,TP135D0 ,TP127D0 ,TP119D0 ,TP142D3 ;
  input TP134D3 ,TP126D3 ,TP118D3 ,TP142D2 ,TP134D2 ,TP126D2 ,TP118D2 ,TP142D1 ,TP134D1 ;
  input TP126D1 ,TP118D1 ,TP142D0 ,TP134D0 ,TP126D0 ,TP118D0 ,TP141D3 ,TP133D3 ,TP125D3 ;
  input TP117D3 ,TP109D3 ,TP141D2 ,TP133D2 ,TP125D2 ,TP117D2 ,TP109D2 ,TP141D1 ,TP133D1 ;
  input TP125D1 ,TP117D1 ,TP109D1 ,TP141D0 ,TP133D0 ,TP125D0 ,TP117D0 ,TP109D0 ,TP140D3 ;
  input TP132D3 ,TP124D3 ,TP116D3 ,TP108D3 ,TP140D2 ,TP132D2 ,TP124D2 ,TP116D2 ,TP108D2 ;
  input TP140D1 ,TP132D1 ,TP124D1 ,TP116D1 ,TP108D1 ,TP140D0 ,TP132D0 ,TP124D0 ,TP116D0 ;
  input TP108D0 ,TP139D3 ,TP139D2 ,TP139D1 ,TP139D0 ,TP138D3 ,TP138D2 ,TP138D1 ,TP138D0 ;
  input TP137D3 ,TP129D3 ,TP137D2 ,TP129D2 ,TP137D1 ,TP129D1 ,TP137D0 ,TP129D0 ,TP131D3 ;
  input TP123D3 ,TP115D3 ,TP107D3 ,TP131D2 ,TP123D2 ,TP115D2 ,TP107D2 ,TP131D1 ,TP123D1 ;
  input TP115D1 ,TP107D1 ,TP131D0 ,TP123D0 ,TP115D0 ,TP107D0 ,TP130D3 ,TP122D3 ,TP114D3 ;
  input TP106D3 ,TP130D2 ,TP122D2 ,TP114D2 ,TP106D2 ,TP130D1 ,TP122D1 ,TP114D1 ,TP106D1 ;
  input TP130D0 ,TP122D0 ,TP114D0 ,TP106D0 ,TP121D3 ,TP113D3 ,TP105D3 ,TP121D2 ,TP113D2 ;
  input TP105D2 ,TP121D1 ,TP113D1 ,TP105D1 ,TP121D0 ,TP113D0 ,TP105D0 ,TP120D3 ,TP112D3 ;
  input TP104D3 ,TP120D2 ,TP112D2 ,TP104D2 ,TP120D1 ,TP112D1 ,TP104D1 ,TP120D0 ,TP112D0 ;
  input TP104D0 ,TP111D3 ,TP103D3 ,TP111D2 ,TP103D2 ,TP111D1 ,TP103D1 ,TP111D0 ,TP103D0 ;
  input TP110D3 ,TP102D3 ,TP110D2 ,TP102D2 ,TP110D1 ,TP102D1 ,TP110D0 ,TP102D0 ,TP101D3 ;
  input TP101D2 ,TP101D1 ,TP101D0 ,TP100D3 ,TP100D2 ,TP100D1 ,TP100D0 ,TP99D3 ,TP99D2 ;
  input TP99D1 ,TP99D0 ,TP98D3 ,TP98D2 ,TP98D1 ,TP98D0 ,TP97D3 ,TP89D3 ,TP97D2 ;
  input TP89D2 ,TP97D1 ,TP89D1 ,TP97D0 ,TP89D0 ,TP96D3 ,TP88D3 ,TP96D2 ,TP88D2 ;
  input TP96D1 ,TP88D1 ,TP96D0 ,TP88D0 ,TP95D3 ,TP87D3 ,TP79D3 ,TP95D2 ,TP87D2 ;
  input TP79D2 ,TP95D1 ,TP87D1 ,TP79D1 ,TP95D0 ,TP87D0 ,TP79D0 ,TP94D3 ,TP86D3 ;
  input TP78D3 ,TP94D2 ,TP86D2 ,TP78D2 ,TP94D1 ,TP86D1 ,TP78D1 ,TP94D0 ,TP86D0 ;
  input TP78D0 ,TP93D3 ,TP85D3 ,TP77D3 ,TP69D3 ,TP93D2 ,TP85D2 ,TP77D2 ,TP69D2 ;
  input TP93D1 ,TP85D1 ,TP77D1 ,TP69D1 ,TP93D0 ,TP85D0 ,TP77D0 ,TP69D0 ,TP92D3 ;
  input TP84D3 ,TP76D3 ,TP68D3 ,TP92D2 ,TP84D2 ,TP76D2 ,TP68D2 ,TP92D1 ,TP84D1 ;
  input TP76D1 ,TP68D1 ,TP92D0 ,TP84D0 ,TP76D0 ,TP68D0 ,TP91D3 ,TP83D3 ,TP75D3 ;
  input TP67D3 ,TP59D3 ,TP91D2 ,TP83D2 ,TP75D2 ,TP67D2 ,TP59D2 ,TP91D1 ,TP83D1 ;
  input TP75D1 ,TP67D1 ,TP59D1 ,TP91D0 ,TP83D0 ,TP75D0 ,TP67D0 ,TP59D0 ,TP90D3 ;
  input TP82D3 ,TP74D3 ,TP66D3 ,TP58D3 ,TP90D2 ,TP82D2 ,TP74D2 ,TP66D2 ,TP58D2 ;
  input TP90D1 ,TP82D1 ,TP74D1 ,TP66D1 ,TP58D1 ,TP90D0 ,TP82D0 ,TP74D0 ,TP66D0 ;
  input TP58D0 ,TP81D3 ,TP73D3 ,TP65D3 ,TP57D3 ,TP49D3 ,TP81D2 ,TP73D2 ,TP65D2 ;
  input TP57D2 ,TP49D2 ,TP81D1 ,TP73D1 ,TP65D1 ,TP57D1 ,TP49D1 ,TP81D0 ,TP73D0 ;
  input TP65D0 ,TP57D0 ,TP49D0 ,TP80D3 ,TP72D3 ,TP64D3 ,TP56D3 ,TP48D3 ,TP80D2 ;
  input TP72D2 ,TP64D2 ,TP56D2 ,TP48D2 ,TP80D1 ,TP72D1 ,TP64D1 ,TP56D1 ,TP48D1 ;
  input TP80D0 ,TP72D0 ,TP64D0 ,TP56D0 ,TP48D0 ,TP71D3 ,TP63D3 ,TP55D3 ,TP47D3 ;
  input TP39D3 ,TP71D2 ,TP63D2 ,TP55D2 ,TP47D2 ,TP39D2 ,TP71D1 ,TP63D1 ,TP55D1 ;
  input TP47D1 ,TP39D1 ,TP71D0 ,TP63D0 ,TP55D0 ,TP47D0 ,TP39D0 ,TP70D3 ,TP62D3 ;
  input TP54D3 ,TP46D3 ,TP38D3 ,TP70D2 ,TP62D2 ,TP54D2 ,TP46D2 ,TP38D2 ,TP70D1 ;
  input TP62D1 ,TP54D1 ,TP46D1 ,TP38D1 ,TP70D0 ,TP62D0 ,TP54D0 ,TP46D0 ,TP38D0 ;
  input TP61D3 ,TP53D3 ,TP45D3 ,TP37D3 ,TP29D3 ,TP61D2 ,TP53D2 ,TP45D2 ,TP37D2 ;
  input TP29D2 ,TP61D1 ,TP53D1 ,TP45D1 ,TP37D1 ,TP29D1 ,TP61D0 ,TP53D0 ,TP45D0 ;
  input TP37D0 ,TP29D0 ,TP60D3 ,TP52D3 ,TP44D3 ,TP36D3 ,TP28D3 ,TP60D2 ,TP52D2 ;
  input TP44D2 ,TP36D2 ,TP28D2 ,TP60D1 ,TP52D1 ,TP44D1 ,TP36D1 ,TP28D1 ,TP60D0 ;
  input TP52D0 ,TP44D0 ,TP36D0 ,TP28D0 ,TP51D3 ,TP43D3 ,TP35D3 ,TP27D3 ,TP19D3 ;
  input TP51D2 ,TP43D2 ,TP35D2 ,TP27D2 ,TP19D2 ,TP51D1 ,TP43D1 ,TP35D1 ,TP27D1 ;
  input TP19D1 ,TP51D0 ,TP43D0 ,TP35D0 ,TP27D0 ,TP19D0 ,TP50D3 ,TP42D3 ,TP34D3 ;
  input TP26D3 ,TP18D3 ,TP50D2 ,TP42D2 ,TP34D2 ,TP26D2 ,TP18D2 ,TP50D1 ,TP42D1 ;
  input TP34D1 ,TP26D1 ,TP18D1 ,TP50D0 ,TP42D0 ,TP34D0 ,TP26D0 ,TP18D0 ,TP41D3 ;
  input TP33D3 ,TP25D3 ,TP17D3 ,TP41D2 ,TP33D2 ,TP25D2 ,TP17D2 ,TP41D1 ,TP33D1 ;
  input TP25D1 ,TP17D1 ,TP41D0 ,TP33D0 ,TP25D0 ,TP17D0 ,TP40D3 ,TP32D3 ,TP24D3 ;
  input TP16D3 ,TP40D2 ,TP32D2 ,TP24D2 ,TP16D2 ,TP40D1 ,TP32D1 ,TP24D1 ,TP16D1 ;
  input TP40D0 ,TP32D0 ,TP24D0 ,TP16D0 ,TP31D3 ,TP23D3 ,TP15D3 ,TP31D2 ,TP23D2 ;
  input TP15D2 ,TP31D1 ,TP23D1 ,TP15D1 ,TP31D0 ,TP23D0 ,TP15D0 ,TP30D3 ,TP22D3 ;
  input TP14D3 ,TP30D2 ,TP22D2 ,TP14D2 ,TP30D1 ,TP22D1 ,TP14D1 ,TP30D0 ,TP22D0 ;
  input TP14D0 ,TP21D3 ,TP13D3 ,TP21D2 ,TP13D2 ,TP21D1 ,TP13D1 ,TP21D0 ,TP13D0 ;
  input TP20D3 ,TP12D3 ,TP20D2 ,TP12D2 ,TP20D1 ,TP12D1 ,TP20D0 ,TP12D0 ,TP11D3 ;
  input TP11D2 ,TP11D1 ,TP11D0 ,TP10D3 ,TP10D2 ,TP10D1 ,TP10D0 ,TP9D3 ,TP9D2 ;
  input TP9D1 ,TP9D0 ,TP8D3 ,TP8D2 ,TP8D1 ,TP8D0 ,TP7D3 ,TP7D2 ,TP7D1 ;
  input TP7D0 ,TP6D3 ,TP6D2 ,TP6D1 ,TP6D0 ,TP5D3 ,TP5D2 ,TP5D1 ,TP5D0 ;
  input TP4D3 ,TP4D2 ,TP4D1 ,TP4D0 ,TP3D3 ,TP3D2 ,TP3D1 ,TP3D0 ,TP2D3 ;
  input TP2D2 ,TP2D1 ,TP2D0 ,TP1D3 ,TP1D2 ,TP1D1 ,TP1D0 ,CLK30MHZ ,BTFLG ;
  input TMSPMD ,TMBTSEL ,RESB ,USBCLK ,USBRD_B ,USBWR0_B ,USBA21 ,USBA20 ,USBA19 ;
  input USBA4 ,USBA3 ,USBA2 ,ICESYSRES_B ,ICECPURES_B ,RESET_B ,EVAOSCMCLK ,EVAOSCRCLK1 ,EVAOSCRCLK2 ;
  input EVAOSCRCLK3 ,TCCONNECT_B ,EACONNECT_B ,TVDDON ,DCE0 ,DCLKSEL1 ,DCER ,DSER ,DWWR ;
  input DWED ,DMRG00 ,DMRG01 ,DMRG10 ,DMRG11 ,DMRG12 ,DREAD ,AF19 ,AF18 ;
  input AF17 ,DA13 ,AF16 ,DA12 ,AF15 ,DA11 ,AF14 ,DA10 ,AF13 ;
  input AF12 ,AF11 ,AF10 ,AF9 ,DA7 ,AF8 ,DA6 ,AF5 ,DA3 ;
  input AF4 ,DA2 ,AF3 ,DA1 ,AF2 ,DA0 ,AF1 ,AF0 ,DRDCLK ;
  input DRDCLKC1 ,DA9 ,DA8 ,SLDFLASH ,LOCK240FAIL ,CLK240M ,CLK120M ;


  output CLK30MHZ_GB ,ICEWAITMEM ,ICENOECC ,ICEFLERR ,RO137 ,RO129 ,RO136 ,RO128 ,RO135 ;
  output RO127 ,RO119 ,RO134 ,RO126 ,RO118 ,RO133 ,RO125 ,RO117 ,RO037 ;
  output RO029 ,RO132 ,RO124 ,RO116 ,RO036 ,RO028 ,RO131 ,RO123 ,RO115 ;
  output RO035 ,RO027 ,RO019 ,RO130 ,RO122 ,RO114 ,RO034 ,RO026 ,RO018 ;
  output RO121 ,RO113 ,RO033 ,RO025 ,RO017 ,RO120 ,RO112 ,RO032 ,RO024 ;
  output RO016 ,RO111 ,RO031 ,RO023 ,RO015 ,RO110 ,RO030 ,RO022 ,RO014 ;
  output RO19 ,RO18 ,RO17 ,RO09 ,RO16 ,RO08 ,RO15 ,RO07 ,RO14 ;
  output RO06 ,RO13 ,RO05 ,RO12 ,RO04 ,RO11 ,RO03 ,RO10 ,RO02 ;
  output RO021 ,RO013 ,RO020 ,RO012 ,RO011 ,RO010 ,RO01 ,RO00 ,WAITFL2 ;
  output TMEMA14 ,CPUPID31 ,CPUPID23 ,CPUPID15 ,CPUPID30 ,CPUPID22 ,CPUPID14 ,CPUPID29 ,CPUPID28 ;
  output CPUPID27 ,CPUPID19 ,CPUPID26 ,CPUPID18 ,CPUPID25 ,CPUPID17 ,CPUPID24 ,CPUPID16 ,CPUPID21 ;
  output CPUPID13 ,CPUPID20 ,CPUPID12 ,CPUPID11 ,CPUPID10 ,CPUPID9 ,CPUPID8 ,CPUPID7 ,CPUPID6 ;
  output CPUPID5 ,CPUPID4 ,CPUPID3 ,CPUPID2 ,CPUPID1 ,CPUPID0 ,ICEIFA31 ,ICEIFA23 ,ICEIFA15 ;
  output ICEIFA30 ,ICEIFA22 ,ICEIFA14 ,ICEIFA29 ,ICEIFA28 ,ICEIFA27 ,ICEIFA19 ,ICEIFA26 ,ICEIFA18 ;
  output ICEIFA25 ,ICEIFA17 ,ICEIFA24 ,ICEIFA16 ,ICEIFA21 ,ICEIFA13 ,ICEIFA20 ,ICEIFA12 ,ICEIFA11 ;
  output ICEIFA10 ,ICEIFA9 ,ICEIFA8 ,ICEIFA7 ,ICEIFA6 ,ICEIFA5 ,ICEIFA4 ,ICEIFA3 ,ICEIFA2 ;
  output ICEIFA1 ,ICEIFA0 ,ICEDI31 ,ICEDI23 ,ICEDI15 ,ICEDI30 ,ICEDI22 ,ICEDI14 ,ICEDI29 ;
  output ICEDI28 ,ICEDI27 ,ICEDI19 ,ICEDI26 ,ICEDI18 ,ICEDI25 ,ICEDI17 ,ICEDI24 ,ICEDI16 ;
  output ICEDI21 ,ICEDI13 ,ICEDI20 ,ICEDI12 ,ICEDI11 ,ICEDI10 ,ICEDI9 ,ICEDI8 ,ICEDI7 ;
  output ICEDI6 ,ICEDI5 ,ICEDI4 ,ICEDI3 ,ICEDI2 ,ICEDI1 ,ICEDI0 ,ICEWR ,VDDLEV7 ;
  output VDDLEV6 ,VDDLEV5 ,VDDLEV4 ,VDDLEV3 ,VDDLEV2 ,VDDLEV1 ,VDDLEV0 ,USBIFWR ,ICECSGREGU ;
  output POCRESB ,TARRESB ,CLK60MHZ ,CLK60MHZLOCK ,CPUMCLK ,CPUSCLK ,CPURCLK1 ,CPURCLK2 ,CPURCLK3 ;
  output STBRELESV ,SVI ,SVMODI ,SVMODIPERI1 ,SVMODIPERI2 ,SVVCOUT7 ,SVVCOUT6 ,SVVCOUT5 ,SVVCOUT4 ;
  output SVVCOUT3 ,SVVCOUT2 ,SVVCOUT1 ,SVVCOUT0 ,SVMODOPBRK ,FLSIZE3 ,FLSIZE2 ,FLSIZE1 ,FLSIZE0 ;
  output RAMSIZE7 ,RAMSIZE6 ,RAMSIZE5 ,RAMSIZE4 ,RAMSIZE3 ,RAMSIZE2 ,RAMSIZE1 ,RAMSIZE0 ,BFSIZE3 ;
  output BFSIZE2 ,BFSIZE1 ,BFSIZE0 ,BMSIZE3 ,BMSIZE2 ,BMSIZE1 ,BMSIZE0 ,DFSIZE1 ,DFSIZE0 ;
  output SELRAMMA ,SELDFADMA ,PSEUDOON31 ,PSEUDOON23 ,PSEUDOON15 ,PSEUDOON30 ,PSEUDOON22 ,PSEUDOON14 ,PSEUDOON29 ;
  output PSEUDOON28 ,PSEUDOON27 ,PSEUDOON19 ,PSEUDOON26 ,PSEUDOON18 ,PSEUDOON25 ,PSEUDOON17 ,PSEUDOON24 ,PSEUDOON16 ;
  output PSEUDOON21 ,PSEUDOON13 ,PSEUDOON20 ,PSEUDOON12 ,PSEUDOON11 ,PSEUDOON10 ,PSEUDOON9 ,PSEUDOON8 ,PSEUDOON7 ;
  output PSEUDOON6 ,PSEUDOON5 ,PSEUDOON4 ,PSEUDOON3 ,PSEUDOON2 ,PSEUDOON1 ,PSEUDOON0 ,PSEUDOANI09 ,PSEUDOANI17 ;
  output PSEUDOANI08 ,PSEUDOANI16 ,PSEUDOANI07 ,PSEUDOANI15 ,PSEUDOANI06 ,PSEUDOANI14 ,PSEUDOANI05 ,PSEUDOANI13 ,PSEUDOANI04 ;
  output PSEUDOANI12 ,PSEUDOANI03 ,PSEUDOANI11 ,PSEUDOANI02 ,PSEUDOANI10 ,PSEUDOANI01 ,PSEUDOANI00 ,PSEUDOANI19 ,PSEUDOANI18 ;
  output ICEMSKDBG ,ICEMSKWAIT ,ICEMSKNMI ,ICEMSKTRAP ,ICEMSKWDT ,ICEMSKLVI ,ICEMSKRETRY ,MDR_RAM15 ,MDR_RAM14 ;
  output MDR_RAM13 ,MDR_RAM12 ,MDR_RAM11 ,MDR_RAM10 ,MDR_RAM9 ,MDR_RAM8 ,MDR_RAM7 ,MDR_RAM6 ,MDR_RAM5 ;
  output MDR_RAM4 ,MDR_RAM3 ,MDR_RAM2 ,MDR_RAM1 ,MDR_RAM0 ,SYSRSOUTB ,PONRESB ,ADDRTD144 ,ADDRTD136 ;
  output ADDRTD128 ,ADDRTD143 ,ADDRTD135 ,ADDRTD127 ,ADDRTD119 ,ADDRTD142 ,ADDRTD134 ,ADDRTD126 ,ADDRTD118 ;
  output ADDRTD141 ,ADDRTD133 ,ADDRTD125 ,ADDRTD117 ,ADDRTD109 ,ADDRTD140 ,ADDRTD132 ,ADDRTD124 ,ADDRTD116 ;
  output ADDRTD108 ,ADDRTD139 ,ADDRTD138 ,ADDRTD137 ,ADDRTD129 ,ADDRTD131 ,ADDRTD123 ,ADDRTD115 ,ADDRTD107 ;
  output ADDRTD130 ,ADDRTD122 ,ADDRTD114 ,ADDRTD106 ,ADDRTD121 ,ADDRTD113 ,ADDRTD105 ,ADDRTD120 ,ADDRTD112 ;
  output ADDRTD104 ,ADDRTD111 ,ADDRTD103 ,ADDRTD110 ,ADDRTD102 ,ADDRTD101 ,ADDRTD100 ,ADDRTD99 ,ADDRTD98 ;
  output ADDRTD97 ,ADDRTD89 ,ADDRTD96 ,ADDRTD88 ,ADDRTD95 ,ADDRTD87 ,ADDRTD79 ,ADDRTD94 ,ADDRTD86 ;
  output ADDRTD78 ,ADDRTD93 ,ADDRTD85 ,ADDRTD77 ,ADDRTD69 ,ADDRTD92 ,ADDRTD84 ,ADDRTD76 ,ADDRTD68 ;
  output ADDRTD91 ,ADDRTD83 ,ADDRTD75 ,ADDRTD67 ,ADDRTD59 ,ADDRTD90 ,ADDRTD82 ,ADDRTD74 ,ADDRTD66 ;
  output ADDRTD58 ,ADDRTD81 ,ADDRTD73 ,ADDRTD65 ,ADDRTD57 ,ADDRTD49 ,ADDRTD80 ,ADDRTD72 ,ADDRTD64 ;
  output ADDRTD56 ,ADDRTD48 ,ADDRTD71 ,ADDRTD63 ,ADDRTD55 ,ADDRTD47 ,ADDRTD39 ,ADDRTD70 ,ADDRTD62 ;
  output ADDRTD54 ,ADDRTD46 ,ADDRTD38 ,ADDRTD61 ,ADDRTD53 ,ADDRTD45 ,ADDRTD37 ,ADDRTD29 ,ADDRTD60 ;
  output ADDRTD52 ,ADDRTD44 ,ADDRTD36 ,ADDRTD28 ,ADDRTD51 ,ADDRTD43 ,ADDRTD35 ,ADDRTD27 ,ADDRTD19 ;
  output ADDRTD50 ,ADDRTD42 ,ADDRTD34 ,ADDRTD26 ,ADDRTD18 ,ADDRTD41 ,ADDRTD33 ,ADDRTD25 ,ADDRTD17 ;
  output ADDRTD40 ,ADDRTD32 ,ADDRTD24 ,ADDRTD16 ,ADDRTD31 ,ADDRTD23 ,ADDRTD15 ,ADDRTD30 ,ADDRTD22 ;
  output ADDRTD14 ,ADDRTD21 ,ADDRTD13 ,ADDRTD20 ,ADDRTD12 ,ADDRTD11 ,ADDRTD10 ,ADDRTD9 ,ADDRTD8 ;
  output ADDRTD7 ,ADDRTD6 ,ADDRTD5 ,ADDRTD4 ,ADDRTD3 ,ADDRTD2 ,ADDRTD1 ,ADDRPINRD ,ADDRPINMD ;
  output ADDRPINLV ,EROMWRB ,EROMRDB ,EROMCSB ,EROMPA2 ,EROMCLK ,EROMPA17 ,EROMPA16 ,EROMPA15 ;
  output EROMPA14 ,EROMPA13 ,EROMPA12 ,EROMPA11 ,EROMPA10 ,EROMPA9 ,EROMPA8 ,EROMPA7 ,EROMPA6 ;
  output EROMPA5 ,EROMPA4 ,EROMPA3 ,EROMPA1 ,EROMPA0 ,RDCLKP1_OUT ,EXA_OUT ,WWR_OUT ,CER_OUT ;
  output SER_OUT ,EXER_OUT ,MRG00_OUT ,MRG01_OUT ,MRG10_OUT ,MRG11_OUT ,MRG12_OUT ,DIS_OUT ,READ_OUT ;
  output FCLK_OUT ,PROGI_OUT ,BFA_OUT ,ICETMSPMD ,ICETMBTSEL ,USBWAIT_B ,TMEMA16 ,TMEMA15 ,TMEMA13 ;
  output TMEMA12 ,TMEMA11 ,TMEMA10 ,TMEMA9 ,TMEMA8 ,TMEMA7 ,TMEMA6 ,TMEMA5 ,TMEMA4 ;
  output TMEMA3 ,TMEMA2 ,TMEMA1 ,TMEMA0 ,TMEMCS_B ,TMEMRD_B ,TMEMWR_B ,TMEMCLK2 ,TMEMCLK1 ;
  output TMEMCLK0 ,TVDDSEL ,LEDTVDD_B ,LEDCLOCK_B ,LEDRUN_B ,LEDRESET_B ,LEDSTANDBY_B ,LEDWAIT_B ,DRO11 ;
  output DRO10 ,DRO9 ,DRO8 ,DRO7 ,DRO6 ,DRO5 ,DRO4 ,DRO3 ,DRO2 ;
  output DRO1 ,DRO0 ,DDIS_OUT ,DRDCLKP1_OUT ,DWWR_OUT ,DCER_OUT ,DSER_OUT ,DMRG00_OUT ,DMRG01_OUT ;
  output DMRG10_OUT ,DMRG11_OUT ,DMRG12_OUT ,DREAD_OUT ,DFCLK_OUT ;


  inout EROMPD3 ,EROMPD2 ,EROMPD1 ,EROMPD0 ,EROMPD31 ,EROMPD23 ,EROMPD15 ,EROMPD30 ,EROMPD22 ;
  inout EROMPD14 ,EROMPD29 ,EROMPD28 ,EROMPD27 ,EROMPD19 ,EROMPD26 ,EROMPD18 ,EROMPD25 ,EROMPD17 ;
  inout EROMPD24 ,EROMPD16 ,EROMPD21 ,EROMPD13 ,EROMPD20 ,EROMPD12 ,EROMPD11 ,EROMPD10 ,EROMPD9 ;
  inout EROMPD8 ,EROMPD7 ,EROMPD6 ,EROMPD5 ,EROMPD4 ,USBD15 ,USBD14 ,USBD13 ,USBD12 ;
  inout USBD11 ,USBD10 ,USBD9 ,USBD8 ,USBD7 ,USBD6 ,USBD5 ,USBD4 ,USBD3 ;
  inout USBD2 ,USBD1 ,USBD0 ,TMEMD3 ,TMEMD2 ,TMEMD1 ,TMEMD0 ,TMEMD107 ,TMEMD106 ;
  inout TMEMD105 ,TMEMD104 ,TMEMD103 ,TMEMD102 ,TMEMD101 ,TMEMD100 ,TMEMD99 ,TMEMD98 ,TMEMD97 ;
  inout TMEMD89 ,TMEMD96 ,TMEMD88 ,TMEMD95 ,TMEMD87 ,TMEMD79 ,TMEMD94 ,TMEMD86 ,TMEMD78 ;
  inout TMEMD93 ,TMEMD85 ,TMEMD77 ,TMEMD69 ,TMEMD92 ,TMEMD84 ,TMEMD76 ,TMEMD68 ,TMEMD91 ;
  inout TMEMD83 ,TMEMD75 ,TMEMD67 ,TMEMD59 ,TMEMD90 ,TMEMD82 ,TMEMD74 ,TMEMD66 ,TMEMD58 ;
  inout TMEMD81 ,TMEMD73 ,TMEMD65 ,TMEMD57 ,TMEMD49 ,TMEMD80 ,TMEMD72 ,TMEMD64 ,TMEMD56 ;
  inout TMEMD48 ,TMEMD71 ,TMEMD63 ,TMEMD55 ,TMEMD47 ,TMEMD39 ,TMEMD70 ,TMEMD62 ,TMEMD54 ;
  inout TMEMD46 ,TMEMD38 ,TMEMD61 ,TMEMD53 ,TMEMD45 ,TMEMD37 ,TMEMD29 ,TMEMD60 ,TMEMD52 ;
  inout TMEMD44 ,TMEMD36 ,TMEMD28 ,TMEMD51 ,TMEMD43 ,TMEMD35 ,TMEMD27 ,TMEMD19 ,TMEMD50 ;
  inout TMEMD42 ,TMEMD34 ,TMEMD26 ,TMEMD18 ,TMEMD41 ,TMEMD33 ,TMEMD25 ,TMEMD17 ,TMEMD40 ;
  inout TMEMD32 ,TMEMD24 ,TMEMD16 ,TMEMD31 ,TMEMD23 ,TMEMD15 ,TMEMD30 ,TMEMD22 ,TMEMD14 ;
  inout TMEMD21 ,TMEMD13 ,TMEMD20 ,TMEMD12 ,TMEMD11 ,TMEMD10 ,TMEMD9 ,TMEMD8 ,TMEMD7 ;
  inout TMEMD6 ,TMEMD5 ,TMEMD4 ;


  wire  CLK30MHZ_GB ,A19 ,A18 ,A17 ,A16 ,A15 ,A14 ,A13 ,A12 ;
  wire  A11 ,A10 ,A9 ,A8 ,A7 ,A6 ,A5 ,A4 ,A3 ;
  wire  A2 ,DW37 ,DW29 ,PA13 ,DW36 ,DW28 ,PA12 ,DW35 ,DW27 ;
  wire  DW19 ,PA11 ,DW34 ,DW26 ,DW18 ,PA10 ,DW33 ,DW25 ,DW17 ;
  wire  DDIS ,DW32 ,DW24 ,DW16 ,DW31 ,DW23 ,DW15 ,DW30 ,DW22 ;
  wire  DW14 ,DW21 ,DW13 ,ALT1 ,DW20 ,DW12 ,DW11 ,DW10 ,DW9 ;
  wire  PA5 ,PC1 ,DW8 ,PA4 ,PC0 ,DW7 ,DIS ,PA3 ,DW6 ;
  wire  PA2 ,DW5 ,DW4 ,DW3 ,DW2 ,DW1 ,MA9 ,DW0 ,MA8 ;
  wire  BEU2 ,MA12 ,BEU1 ,MA11 ,BEU0 ,MA10 ,READ ,TAG8 ,MRG00 ;
  wire  TI3D0 ,MRG01 ,TI3D1 ,MRG10 ,TI3D2 ,MRG11 ,TI3D3 ,MRG12 ,TI4D0 ;
  wire  WWR ,CLKSEL1 ,RDCLKP1 ,FCLK ,PA19 ,PC11 ,PROGI ,USBA1 ,CER ;
  wire  MA2 ,SER ,CE0 ,AF6 ,DA4 ,CE1 ,AF7 ,DA5 ,EXA ;
  wire  WED ,EXCH ,MDW0 ,FLMD0 ,FLMA6 ,SELRO1 ,BRSAM ,ICEWAITMEM ,ICENOECC ;
  wire  ICEFLERR ,RO137 ,RO129 ,EXMA3 ,TAG21 ,TAG13 ,RO136 ,RO128 ,EXMA2 ;
  wire  TAG20 ,TAG12 ,RO135 ,RO127 ,RO119 ,EXMA1 ,TAG11 ,RO134 ,RO126 ;
  wire  RO118 ,EXMA0 ,TAG10 ,RO133 ,RO125 ,RO117 ,RO037 ,RO029 ,RO132 ;
  wire  RO124 ,RO116 ,RO036 ,RO028 ,RO131 ,RO123 ,RO115 ,RO035 ,RO027 ;
  wire  RO019 ,RO130 ,RO122 ,RO114 ,RO034 ,RO026 ,RO018 ,RO121 ,RO113 ;
  wire  RO033 ,RO025 ,RO017 ,RO120 ,RO112 ,RO032 ,RO024 ,RO016 ,RO111 ;
  wire  RO031 ,RO023 ,RO015 ,RO110 ,RO030 ,RO022 ,RO014 ,RO19 ,TAG5 ;
  wire  RO18 ,TAG4 ,RO17 ,RO09 ,TAG3 ,RO16 ,RO08 ,TAG2 ,RO15 ;
  wire  RO07 ,TAG1 ,RO14 ,RO06 ,TAG0 ,RO13 ,RO05 ,RO12 ,RO04 ;
  wire  RO11 ,RO03 ,MDW9 ,RO10 ,RO02 ,MDW8 ,RO021 ,RO013 ,RO020 ;
  wire  RO012 ,CPURD ,RO011 ,RO010 ,RO01 ,MDW7 ,RO00 ,MDW6 ,WAITFL2 ;
  wire  SLFLASH ,TMEMA14 ,GDRAMWR ,CIBPID31 ,CIBPID23 ,CIBPID15 ,CIBPID30 ,CIBPID22 ,CIBPID14 ;
  wire  CIBPID29 ,CIBPID28 ,CIBPID27 ,CIBPID19 ,CIBPID26 ,CIBPID18 ,CIBPID25 ,CIBPID17 ,CIBPID24 ;
  wire  CIBPID16 ,CIBPID21 ,CIBPID13 ,CIBPID20 ,CIBPID12 ,CIBPID11 ,CIBPID10 ,CIBPID9 ,CIBPID8 ;
  wire  CIBPID7 ,CIBPID6 ,CIBPID5 ,CIBPID4 ,CIBPID3 ,CIBPID2 ,CIBPID1 ,CIBPID0 ,CPUPID31 ;
  wire  CPUPID23 ,CPUPID15 ,CPUPID30 ,CPUPID22 ,CPUPID14 ,CPUPID29 ,CPUPID28 ,CPUPID27 ,CPUPID19 ;
  wire  CPUPID26 ,CPUPID18 ,CPUPID25 ,CPUPID17 ,CPUPID24 ,CPUPID16 ,CPUPID21 ,CPUPID13 ,CPUPID20 ;
  wire  CPUPID12 ,CPUPID11 ,CPUPID10 ,CPUPID9 ,CPUPID8 ,CPUPID7 ,CPUPID6 ,CPUPID5 ,CPUPID4 ;
  wire  CPUPID3 ,CPUPID2 ,CPUPID1 ,CPUMASK ,CPUPID0 ,EMEMRAMCLK ,ICEIFA31 ,ICEIFA23 ,ICEIFA15 ;
  wire  ICEDOD11 ,ICEDOB27 ,ICEDOB19 ,ICEDOC31 ,ICEDOC23 ,ICEDOC15 ,ICEIFA30 ,ICEIFA22 ,ICEIFA14 ;
  wire  ICEDOD10 ,ICEDOB26 ,ICEDOB18 ,ICEDOC30 ,ICEDOC22 ,ICEDOC14 ,ICEIFA29 ,ICEDOE21 ,ICEDOE13 ;
  wire  ICEDOD25 ,ICEDOD17 ,ICEDOC29 ,ICEIFA28 ,ICEDOE20 ,ICEDOE12 ,ICEDOD24 ,ICEDOD16 ,ICEDOC28 ;
  wire  ICEIFA27 ,ICEIFA19 ,ICEDOE11 ,ICEDOD31 ,ICEDOD23 ,ICEDOD15 ,ICEDOC27 ,ICEDOC19 ,ICEIFA26 ;
  wire  ICEIFA18 ,ICEDOE10 ,ICEDOD30 ,ICEDOD22 ,ICEDOD14 ,ICEDOC26 ,ICEDOC18 ,ICEIFA25 ,ICEIFA17 ;
  wire  ICEDOD21 ,ICEDOD13 ,ICEDOB29 ,ICEDOC25 ,ICEDOC17 ,ICEIFA24 ,ICEIFA16 ,ICEDOD20 ,ICEDOD12 ;
  wire  ICEDOB28 ,ICEDOC24 ,ICEDOC16 ,ICEIFA21 ,ICEIFA13 ,ICEDOA29 ,ICEDOB25 ,ICEDOB17 ,ICEDOC21 ;
  wire  ICEDOC13 ,ICEIFA20 ,ICEIFA12 ,ICEDOA28 ,ICEDOB24 ,ICEDOB16 ,ICEDOC20 ,ICEDOC12 ,ICEIFA11 ;
  wire  ICEDOA27 ,ICEDOA19 ,ICEDOB31 ,ICEDOB23 ,ICEDOB15 ,ICEDOC11 ,ICEIFA10 ,ICEDOA26 ,ICEDOA18 ;
  wire  ICEDOB30 ,ICEDOB22 ,ICEDOB14 ,ICEDOC10 ,ICEIFA9 ,ICEDOE5 ,ICEDOD7 ,ICEDOC9 ,ICEDOF3 ;
  wire  ICEDOG1 ,ICEIFA8 ,ICEDOE4 ,ICEDOD6 ,ICEDOC8 ,ICEDOF2 ,ICEDOG0 ,ICEIFA7 ,ICEDOE3 ;
  wire  ICEDOD5 ,ICEDOB9 ,ICEDOC7 ,ICEDOF1 ,ICEIFA6 ,ICEDOE2 ,ICEDOD4 ,ICEDOB8 ,ICEDOC6 ;
  wire  ICEDOF0 ,ICEIFA5 ,ICEDOA9 ,ICEDOE1 ,ICEDOD3 ,ICEDOB7 ,ICEDOC5 ,ICEIFA4 ,ICEDOA8 ;
  wire  ICEDOE0 ,ICEDOD2 ,ICEDOB6 ,ICEDOC4 ,ICEIFA3 ,ICEDOA7 ,ICEDOD1 ,ICEDOB5 ,ICEDOC3 ;
  wire  ICEIFA2 ,ICEDOA6 ,ICEDOD0 ,ICEDOB4 ,ICEDOC2 ,ICEIFA1 ,ICEDOA5 ,ICEDOB3 ,ICEDOC1 ;
  wire  ICEIFA0 ,ICEDOA4 ,ICEDOB2 ,ICEDOC0 ,ICEDI31 ,ICEDI23 ,ICEDI15 ,IDADR11 ,ICEDI30 ;
  wire  ICEDI22 ,ICEDI14 ,IDADR10 ,ICEDI29 ,IDADR25 ,IDADR17 ,ICEDI28 ,IDADR24 ,IDADR16 ;
  wire  ICEDI27 ,ICEDI19 ,IDADR31 ,IDADR23 ,IDADR15 ,ICEDI26 ,ICEDI18 ,IDADR30 ,IDADR22 ;
  wire  IDADR14 ,ICEDI25 ,ICEDI17 ,IDADR21 ,IDADR13 ,ICEDI24 ,ICEDI16 ,IDADR20 ,IDADR12 ;
  wire  ICEDI21 ,ICEDI13 ,ICEDI20 ,ICEDI12 ,ICEDI11 ,ICEDI10 ,ICEDI9 ,IDADR7 ,ICEDI8 ;
  wire  IDADR6 ,ICEDI7 ,IDADR5 ,ICEDI6 ,IDADR4 ,ICEDI5 ,IDADR3 ,ICEDI4 ,IDADR2 ;
  wire  ICEDI3 ,IDADR1 ,ICEDI2 ,IDADR0 ,ICEDI1 ,ICEDI0 ,ICEWR ,ICEDOP31 ,ICEDOP23 ;
  wire  ICEDOP15 ,ICEDOQ11 ,ICEDOP30 ,ICEDOP22 ,ICEDOP14 ,ICEDOQ10 ,ICEDOP29 ,ICEDOQ25 ,ICEDOQ17 ;
  wire  ICEDOR21 ,ICEDOR13 ,ICEDOP28 ,ICEDOQ24 ,ICEDOQ16 ,ICEDOR20 ,ICEDOR12 ,ICEDOP27 ,ICEDOP19 ;
  wire  ICEDOQ31 ,ICEDOQ23 ,ICEDOQ15 ,ICEDOR11 ,ICEDOP26 ,ICEDOP18 ,ICEDOQ30 ,ICEDOQ22 ,ICEDOQ14 ;
  wire  ICEDOR10 ,ICEDOP25 ,ICEDOP17 ,ICEDOQ21 ,ICEDOQ13 ,ICEDOP24 ,ICEDOP16 ,ICEDOQ20 ,ICEDOQ12 ;
  wire  ICEDOP21 ,ICEDOP13 ,ICEDON29 ,ICEDOP20 ,ICEDOP12 ,ICEDON28 ,ICEDOP11 ,ICEDON27 ,ICEDON19 ;
  wire  ICEDOP10 ,ICEDON26 ,ICEDON18 ,ICEDOP9 ,ICEDOQ7 ,ICEDOS3 ,ICEDOT1 ,ICEDOR5 ,ICEDOP8 ;
  wire  ICEDOQ6 ,ICEDOS2 ,ICEDOT0 ,ICEDOR4 ,ICEDOP7 ,ICEDOQ5 ,ICEDOS1 ,ICEDOR3 ,ICEDOP6 ;
  wire  ICEDOQ4 ,ICEDOS0 ,ICEDOR2 ,ICEDOP5 ,ICEDOQ3 ,ICEDON9 ,ICEDOR1 ,ICEDOP4 ,ICEDOQ2 ;
  wire  ICEDON8 ,ICEDOR0 ,ICEDOP3 ,ICEDOQ1 ,ICEDON7 ,ICEDOM9 ,ICEDOP2 ,ICEDOQ0 ,ICEDON6 ;
  wire  ICEDOM8 ,ICEDOP1 ,ICEDON5 ,ICEDOM7 ,ICEDOL9 ,ICEDOP0 ,ICEDON4 ,ICEDOM6 ,ICEDOL8 ;
  wire  ICEDOA31 ,ICEDOA23 ,ICEDOA15 ,ICEDOB11 ,ICEDOA30 ,ICEDOA22 ,ICEDOA14 ,ICEDOB10 ,ICEDOA25 ;
  wire  ICEDOA17 ,ICEDOB21 ,ICEDOB13 ,ICEDOA24 ,ICEDOA16 ,ICEDOB20 ,ICEDOB12 ,ICEDOA21 ,ICEDOA13 ;
  wire  ICEDOA20 ,ICEDOA12 ,ICEDOA11 ,ICEDOA10 ,ICEDOA3 ,ICEDOB1 ,ICEDOA2 ,ICEDOB0 ,ICEDOA1 ;
  wire  ICEDOA0 ,VDDLEV7 ,VDDLEV6 ,VDDLEV5 ,VDDLEV4 ,VDDLEV3 ,VDDLEV2 ,VDDLEV1 ,VDDLEV0 ;
  wire  USBIFWR ,ICECSGREGU ,POCRESB ,TARRESB ,CPUPRCLK2 ,CPUTMCLK ,CPUTSCLK ,CPURCLK1SEL ,CLK60MHZ ;
  wire  CLK60MHZLOCK ,CPUMCLK ,CPUSCLK ,CPURCLK1 ,CPURCLK2 ,CPURCLK3 ,SOFTBRK ,SVINTACK ,STBRELESV ;
  wire  SVI ,SVMODI ,SVMODIPERI1 ,SVMODIPERI2 ,SVVCOUT7 ,SVVCOUT6 ,SVVCOUT5 ,SVVCOUT4 ,SVVCOUT3 ;
  wire  SVVCOUT2 ,SVVCOUT1 ,SVVCOUT0 ,SVMODOPBRK ,IDADR29 ,IDADR28 ,IDADR27 ,IDADR19 ,IDADR26 ;
  wire  IDADR18 ,IDADR9 ,IDADR8 ,PERISVIB ,FLSIZE3 ,FLSIZE2 ,FLSIZE1 ,FLSIZE0 ,RAMSIZE7 ;
  wire  RAMSIZE6 ,RAMSIZE5 ,RAMSIZE4 ,RAMSIZE3 ,RAMSIZE2 ,RAMSIZE1 ,RAMSIZE0 ,BFSIZE3 ,BFSIZE2 ;
  wire  BFSIZE1 ,BFSIZE0 ,BMSIZE3 ,BRKMDR1 ,BMSIZE2 ,BRKMDR0 ,BMSIZE1 ,BMSIZE0 ,DFSIZE1 ;
  wire  DFSIZE0 ,SELRAMMA ,SELDFADMA ,PSEUDOON31 ,PSEUDOON23 ,PSEUDOON15 ,PSEUDOON30 ,PSEUDOON22 ,PSEUDOON14 ;
  wire  PSEUDOON29 ,PSEUDOON28 ,PSEUDOON27 ,PSEUDOON19 ,PSEUDOON26 ,PSEUDOON18 ,PSEUDOON25 ,PSEUDOON17 ,PSEUDOON24 ;
  wire  PSEUDOON16 ,PSEUDOON21 ,PSEUDOON13 ,PSEUDOON20 ,PSEUDOON12 ,PSEUDOON11 ,PSEUDOON10 ,PSEUDOON9 ,PSEUDOON8 ;
  wire  PSEUDOON7 ,PSEUDOON6 ,PSEUDOON5 ,PSEUDOON4 ,PSEUDOON3 ,PSEUDOON2 ,PSEUDOON1 ,PSEUDOON0 ,PSEUDOANI09 ;
  wire  PSEUDOANI17 ,PSEUDOANI08 ,PSEUDOANI16 ,PSEUDOANI07 ,PSEUDOANI15 ,PSEUDOANI06 ,PSEUDOANI14 ,PSEUDOANI05 ,PSEUDOANI13 ;
  wire  PSEUDOANI04 ,PSEUDOANI12 ,PSEUDOANI03 ,PSEUDOANI11 ,PSEUDOANI02 ,PSEUDOANI10 ,PSEUDOANI01 ,PSEUDOANI00 ,PSEUDOANI19 ;
  wire  PSEUDOANI18 ,ICEMSKDBG ,ICEMSKWAIT ,ICEMSKNMI ,ICEMSKTRAP ,ICEMSKWDT ,ICEMSKLVI ,ICEMSKRETRY ,MDR_RAM15 ;
  wire  MDR_RAM14 ,MDR_RAM13 ,MDR_RAM12 ,MDR_RAM11 ,MDR_RAM10 ,MDR_RAM9 ,MDR_RAM8 ,MDR_RAM7 ,MDR_RAM6 ;
  wire  MDR_RAM5 ,MDR_RAM4 ,MDR_RAM3 ,MDR_RAM2 ,MDR_RAM1 ,MDR_RAM0 ,CPUWR ,TI1D0 ,WDOP ;
  wire  SVMOD ,SVMODF ,STAGEADR1 ,STAGEADR0 ,PCWAITF ,SKIPEXE ,FCHRAM ,FLREAD ,IMDR10 ;
  wire  FLREADB3 ,FLREADB2 ,FLREADB1 ,FLREADB0 ,CPURSOUTB ,BASECK ,PREFIX ,WAITEXM ,OCDWAIT ;
  wire  MEMMDR6 ,BRAMEN ,BFA ,BFAEN ,INTACK ,DMAACK ,DFMDR1 ,SLEXM ,IDPOP ;
  wire  MDW10 ,IMDR2 ,SPINC ,SPDEC ,SPREL ,CPUMISAL ,SLMEM ,FLSPMD ,STPST ;
  wire  HLTST ,MA15 ,MA14 ,MA13 ,MA7 ,MA6 ,MA5 ,MA4 ,MA3 ;
  wire  MA1 ,MA0 ,MDW15 ,IMDR7 ,MDW14 ,IMDR6 ,MDW13 ,IMDR5 ,MDW12 ;
  wire  IMDR4 ,MDW11 ,IMDR3 ,MDW5 ,MDW4 ,MDW3 ,MDW2 ,DOWN ,MDW1 ;
  wire  PA18 ,PC10 ,PA17 ,PA16 ,PA15 ,PA14 ,PA9 ,PC5 ,PA8 ;
  wire  PC4 ,PA7 ,PC3 ,PA6 ,PC2 ,PC19 ,PC18 ,PC17 ,PC16 ;
  wire  PC15 ,PC14 ,PC13 ,PC12 ,PC9 ,PC8 ,PC7 ,PC6 ,IMDR15 ;
  wire  IMDR14 ,IMDR13 ,IMDR12 ,IMDR11 ,IMDR9 ,IMDR8 ,IMDR1 ,IMDR0 ,SLBMEM ;
  wire  SYSRSOUTB ,PONRESB ,CPUPRCLK3 ,LOCKFAIL5 ,LOCKFAIL6 ,LOCKFAIL7 ,LOCKFAIL8 ,LOCKFAIL9 ,LOCKFAIL10 ;
  wire  LOCKFAIL11 ,LOCKFAIL12 ,LOCKFAIL20 ,LOCKFAIL13 ,LOCKFAIL21 ,LOCKFAIL14 ,LOCKFAIL22 ,LOCKFAIL30 ,LOCKFAIL15 ;
  wire  LOCKFAIL23 ,LOCKFAIL16 ,LOCKFAIL24 ,LOCKFAIL17 ,LOCKFAIL25 ,LOCKFAIL18 ,LOCKFAIL26 ,LOCKFAIL19 ,LOCKFAIL27 ;
  wire  LOCKFAIL28 ,LOCKFAIL29 ,IDVER31 ,IDVER23 ,IDVER15 ,IDVER30 ,IDVER22 ,IDVER14 ,IDVER29 ;
  wire  IDVER28 ,IDVER27 ,IDVER19 ,IDVER26 ,IDVER18 ,IDVER25 ,IDVER17 ,IDVER24 ,IDVER16 ;
  wire  IDVER21 ,IDVER13 ,IDVER20 ,IDVER12 ,IDVER11 ,IDVER10 ,IDVER9 ,IDVER8 ,IDVER7 ;
  wire  IDVER6 ,IDVER5 ,IDVER4 ,IDVER3 ,IDVER2 ,IDVER1 ,IDVER0 ,ADDRTD144 ,ADDRTD136 ;
  wire  ADDRTD128 ,ADDRTD143 ,ADDRTD135 ,ADDRTD127 ,ADDRTD119 ,ADDRTD142 ,ADDRTD134 ,ADDRTD126 ,ADDRTD118 ;
  wire  ADDRTD141 ,ADDRTD133 ,ADDRTD125 ,ADDRTD117 ,ADDRTD109 ,ADDRTD140 ,ADDRTD132 ,ADDRTD124 ,ADDRTD116 ;
  wire  ADDRTD108 ,ADDRTD139 ,ADDRTD138 ,ADDRTD137 ,ADDRTD129 ,ADDRTD131 ,ADDRTD123 ,ADDRTD115 ,ADDRTD107 ;
  wire  ADDRTD130 ,ADDRTD122 ,ADDRTD114 ,ADDRTD106 ,ADDRTD121 ,ADDRTD113 ,ADDRTD105 ,ADDRTD120 ,ADDRTD112 ;
  wire  ADDRTD104 ,ADDRTD111 ,ADDRTD103 ,ADDRTD110 ,ADDRTD102 ,ADDRTD101 ,ADDRTD100 ,ADDRTD99 ,ADDRTD98 ;
  wire  ADDRTD97 ,ADDRTD89 ,ADDRTD96 ,ADDRTD88 ,ADDRTD95 ,ADDRTD87 ,ADDRTD79 ,ADDRTD94 ,ADDRTD86 ;
  wire  ADDRTD78 ,ADDRTD93 ,ADDRTD85 ,ADDRTD77 ,ADDRTD69 ,ADDRTD92 ,ADDRTD84 ,ADDRTD76 ,ADDRTD68 ;
  wire  ADDRTD91 ,ADDRTD83 ,ADDRTD75 ,ADDRTD67 ,ADDRTD59 ,ADDRTD90 ,ADDRTD82 ,ADDRTD74 ,ADDRTD66 ;
  wire  ADDRTD58 ,ADDRTD81 ,ADDRTD73 ,ADDRTD65 ,ADDRTD57 ,ADDRTD49 ,ADDRTD80 ,ADDRTD72 ,ADDRTD64 ;
  wire  ADDRTD56 ,ADDRTD48 ,ADDRTD71 ,ADDRTD63 ,ADDRTD55 ,ADDRTD47 ,ADDRTD39 ,ADDRTD70 ,ADDRTD62 ;
  wire  ADDRTD54 ,ADDRTD46 ,ADDRTD38 ,ADDRTD61 ,ADDRTD53 ,ADDRTD45 ,ADDRTD37 ,ADDRTD29 ,ADDRTD60 ;
  wire  ADDRTD52 ,ADDRTD44 ,ADDRTD36 ,ADDRTD28 ,ADDRTD51 ,ADDRTD43 ,ADDRTD35 ,ADDRTD27 ,ADDRTD19 ;
  wire  ADDRTD50 ,ADDRTD42 ,ADDRTD34 ,ADDRTD26 ,ADDRTD18 ,ADDRTD41 ,ADDRTD33 ,ADDRTD25 ,ADDRTD17 ;
  wire  ADDRTD40 ,ADDRTD32 ,ADDRTD24 ,ADDRTD16 ,ADDRTD31 ,ADDRTD23 ,ADDRTD15 ,ADDRTD30 ,ADDRTD22 ;
  wire  ADDRTD14 ,ADDRTD21 ,ADDRTD13 ,ADDRTD20 ,ADDRTD12 ,ADDRTD11 ,ADDRTD10 ,ADDRTD9 ,ADDRTD8 ;
  wire  ADDRTD7 ,ADDRTD6 ,ADDRTD5 ,ADDRTD4 ,ADDRTD3 ,ADDRTD2 ,ADDRTD1 ,ADDRPINRD ,ADDRPINMD ;
  wire  ADDRPINLV ,TP144D3 ,TP136D3 ,TP128D3 ,TP144D2 ,TP136D2 ,TP128D2 ,TP144D1 ,TP136D1 ;
  wire  TP128D1 ,TP144D0 ,TP136D0 ,TP128D0 ,TP143D3 ,TP135D3 ,TP127D3 ,TP119D3 ,TP143D2 ;
  wire  TP135D2 ,TP127D2 ,TP119D2 ,TP143D1 ,TP135D1 ,TP127D1 ,TP119D1 ,TP143D0 ,TP135D0 ;
  wire  TP127D0 ,TP119D0 ,TP142D3 ,TP134D3 ,TP126D3 ,TP118D3 ,TP142D2 ,TP134D2 ,TP126D2 ;
  wire  TP118D2 ,TP142D1 ,TP134D1 ,TP126D1 ,TP118D1 ,TP142D0 ,TP134D0 ,TP126D0 ,TP118D0 ;
  wire  TP141D3 ,TP133D3 ,TP125D3 ,TP117D3 ,TP109D3 ,TP141D2 ,TP133D2 ,TP125D2 ,TP117D2 ;
  wire  TP109D2 ,TP141D1 ,TP133D1 ,TP125D1 ,TP117D1 ,TP109D1 ,TP141D0 ,TP133D0 ,TP125D0 ;
  wire  TP117D0 ,TP109D0 ,TP140D3 ,TP132D3 ,TP124D3 ,TP116D3 ,TP108D3 ,TP140D2 ,TP132D2 ;
  wire  TP124D2 ,TP116D2 ,TP108D2 ,TP140D1 ,TP132D1 ,TP124D1 ,TP116D1 ,TP108D1 ,TP140D0 ;
  wire  TP132D0 ,TP124D0 ,TP116D0 ,TP108D0 ,TP139D3 ,TP139D2 ,TP139D1 ,TP139D0 ,TP138D3 ;
  wire  TP138D2 ,TP138D1 ,TP138D0 ,TP137D3 ,TP129D3 ,TP137D2 ,TP129D2 ,TP137D1 ,TP129D1 ;
  wire  TP137D0 ,TP129D0 ,ETVDDON ,TP131D3 ,TP123D3 ,TP115D3 ,TP107D3 ,TP131D2 ,TP123D2 ;
  wire  TP115D2 ,TP107D2 ,TP131D1 ,TP123D1 ,TP115D1 ,TP107D1 ,TP131D0 ,TP123D0 ,TP115D0 ;
  wire  TP107D0 ,TP130D3 ,TP122D3 ,TP114D3 ,TP106D3 ,TP130D2 ,TP122D2 ,TP114D2 ,TP106D2 ;
  wire  TP130D1 ,TP122D1 ,TP114D1 ,TP106D1 ,TP130D0 ,TP122D0 ,TP114D0 ,TP106D0 ,TP121D3 ;
  wire  TP113D3 ,TP105D3 ,TP121D2 ,TP113D2 ,TP105D2 ,TP121D1 ,TP113D1 ,TP105D1 ,TP121D0 ;
  wire  TP113D0 ,TP105D0 ,TP120D3 ,TP112D3 ,TP104D3 ,TP120D2 ,TP112D2 ,TP104D2 ,EROMWRB ;
  wire  TP120D1 ,TP112D1 ,TP104D1 ,TP120D0 ,TP112D0 ,TP104D0 ,TP111D3 ,TP103D3 ,TP111D2 ;
  wire  TP103D2 ,TP111D1 ,TP103D1 ,TP111D0 ,TP103D0 ,TP110D3 ,TP102D3 ,TP110D2 ,TP102D2 ;
  wire  TP110D1 ,TP102D1 ,TP110D0 ,TP102D0 ,TP101D3 ,TP101D2 ,TP101D1 ,TP101D0 ,TP100D3 ;
  wire  TP100D2 ,TP100D1 ,TP100D0 ,TP99D3 ,TP99D2 ,TP99D1 ,TP99D0 ,TP98D3 ,TP98D2 ;
  wire  TP98D1 ,TP98D0 ,TP97D3 ,TP89D3 ,TP97D2 ,TP89D2 ,TP97D1 ,TP89D1 ,TP97D0 ;
  wire  TP89D0 ,TP96D3 ,TP88D3 ,TP96D2 ,TP88D2 ,TP96D1 ,TP88D1 ,TP96D0 ,TP88D0 ;
  wire  TP95D3 ,TP87D3 ,TP79D3 ,TP95D2 ,TP87D2 ,TP79D2 ,TP95D1 ,TP87D1 ,TP79D1 ;
  wire  TP95D0 ,TP87D0 ,TP79D0 ,TP94D3 ,TP86D3 ,TP78D3 ,TP94D2 ,TP86D2 ,TP78D2 ;
  wire  TP94D1 ,TP86D1 ,TP78D1 ,TP94D0 ,TP86D0 ,TP78D0 ,TP93D3 ,TP85D3 ,TP77D3 ;
  wire  TP69D3 ,TP93D2 ,TP85D2 ,TP77D2 ,TP69D2 ,TP93D1 ,TP85D1 ,TP77D1 ,TP69D1 ;
  wire  TP93D0 ,TP85D0 ,TP77D0 ,TP69D0 ,TP92D3 ,TP84D3 ,TP76D3 ,TP68D3 ,TP92D2 ;
  wire  TP84D2 ,TP76D2 ,TP68D2 ,TP92D1 ,TP84D1 ,TP76D1 ,TP68D1 ,TP92D0 ,TP84D0 ;
  wire  TP76D0 ,TP68D0 ,TP91D3 ,TP83D3 ,TP75D3 ,TP67D3 ,TP59D3 ,TP91D2 ,TP83D2 ;
  wire  TP75D2 ,TP67D2 ,TP59D2 ,TP91D1 ,TP83D1 ,TP75D1 ,TP67D1 ,TP59D1 ,TP91D0 ;
  wire  TP83D0 ,TP75D0 ,TP67D0 ,TP59D0 ,TP90D3 ,TP82D3 ,TP74D3 ,TP66D3 ,TP58D3 ;
  wire  TP90D2 ,TP82D2 ,TP74D2 ,TP66D2 ,TP58D2 ,TP90D1 ,TP82D1 ,TP74D1 ,TP66D1 ;
  wire  TP58D1 ,TP90D0 ,TP82D0 ,TP74D0 ,TP66D0 ,TP58D0 ,TP81D3 ,TP73D3 ,TP65D3 ;
  wire  TP57D3 ,TP49D3 ,TP81D2 ,TP73D2 ,TP65D2 ,TP57D2 ,TP49D2 ,TP81D1 ,TP73D1 ;
  wire  TP65D1 ,TP57D1 ,TP49D1 ,TP81D0 ,TP73D0 ,TP65D0 ,TP57D0 ,TP49D0 ,TP80D3 ;
  wire  TP72D3 ,TP64D3 ,TP56D3 ,TP48D3 ,TP80D2 ,TP72D2 ,TP64D2 ,TP56D2 ,TP48D2 ;
  wire  TP80D1 ,TP72D1 ,TP64D1 ,TP56D1 ,TP48D1 ,TP80D0 ,TP72D0 ,TP64D0 ,TP56D0 ;
  wire  TP48D0 ,TP71D3 ,TP63D3 ,TP55D3 ,TP47D3 ,TP39D3 ,TP71D2 ,TP63D2 ,TP55D2 ;
  wire  TP47D2 ,TP39D2 ,TP71D1 ,TP63D1 ,TP55D1 ,TP47D1 ,TP39D1 ,TP71D0 ,TP63D0 ;
  wire  TP55D0 ,TP47D0 ,TP39D0 ,TP70D3 ,TP62D3 ,TP54D3 ,TP46D3 ,TP38D3 ,TP70D2 ;
  wire  TP62D2 ,TP54D2 ,TP46D2 ,TP38D2 ,TP70D1 ,TP62D1 ,TP54D1 ,TP46D1 ,TP38D1 ;
  wire  TP70D0 ,TP62D0 ,TP54D0 ,TP46D0 ,TP38D0 ,TP61D3 ,TP53D3 ,TP45D3 ,TP37D3 ;
  wire  TP29D3 ,TP61D2 ,TP53D2 ,TP45D2 ,TP37D2 ,TP29D2 ,TP61D1 ,TP53D1 ,TP45D1 ;
  wire  TP37D1 ,TP29D1 ,TP61D0 ,TP53D0 ,TP45D0 ,TP37D0 ,TP29D0 ,TP60D3 ,TP52D3 ;
  wire  TP44D3 ,TP36D3 ,TP28D3 ,TP60D2 ,TP52D2 ,TP44D2 ,TP36D2 ,TP28D2 ,TP60D1 ;
  wire  TP52D1 ,TP44D1 ,TP36D1 ,TP28D1 ,TP60D0 ,TP52D0 ,TP44D0 ,TP36D0 ,TP28D0 ;
  wire  TP51D3 ,TP43D3 ,TP35D3 ,TP27D3 ,TP19D3 ,TP51D2 ,TP43D2 ,TP35D2 ,TP27D2 ;
  wire  TP19D2 ,TP51D1 ,TP43D1 ,TP35D1 ,TP27D1 ,TP19D1 ,TP51D0 ,TP43D0 ,TP35D0 ;
  wire  TP27D0 ,TP19D0 ,TP50D3 ,TP42D3 ,TP34D3 ,TP26D3 ,TP18D3 ,TP50D2 ,TP42D2 ;
  wire  TP34D2 ,TP26D2 ,TP18D2 ,TP50D1 ,TP42D1 ,TP34D1 ,TP26D1 ,TP18D1 ,TP50D0 ;
  wire  TP42D0 ,TP34D0 ,TP26D0 ,TP18D0 ,TP41D3 ,TP33D3 ,TP25D3 ,TP17D3 ,TP41D2 ;
  wire  TP33D2 ,TP25D2 ,TP17D2 ,TP41D1 ,TP33D1 ,TP25D1 ,TP17D1 ,TP41D0 ,TP33D0 ;
  wire  TP25D0 ,TP17D0 ,TP40D3 ,TP32D3 ,TP24D3 ,TP16D3 ,TP40D2 ,TP32D2 ,TP24D2 ;
  wire  TP16D2 ,TP40D1 ,TP32D1 ,TP24D1 ,TP16D1 ,TP40D0 ,TP32D0 ,TP24D0 ,TP16D0 ;
  wire  TP31D3 ,TP23D3 ,TP15D3 ,TP31D2 ,TP23D2 ,TP15D2 ,TP31D1 ,TP23D1 ,TP15D1 ;
  wire  TP31D0 ,TP23D0 ,TP15D0 ,TP30D3 ,TP22D3 ,TP14D3 ,TP30D2 ,TP22D2 ,TP14D2 ;
  wire  TP30D1 ,TP22D1 ,TP14D1 ,TP30D0 ,TP22D0 ,TP14D0 ,TP21D3 ,TP13D3 ,TP21D2 ;
  wire  TP13D2 ,TP21D1 ,TP13D1 ,TP21D0 ,TP13D0 ,TP20D3 ,TP12D3 ,TP20D2 ,TP12D2 ;
  wire  TP20D1 ,TP12D1 ,TP20D0 ,TP12D0 ,TP11D3 ,TP11D2 ,TP11D1 ,TP11D0 ,TP10D3 ;
  wire  TP10D2 ,TP10D1 ,TP10D0 ,TP9D3 ,TP9D2 ,TP9D1 ,TP9D0 ,TP8D3 ,TP8D2 ;
  wire  TP8D1 ,TP8D0 ,TP7D3 ,TP7D2 ,TP7D1 ,TP7D0 ,TP6D3 ,TP6D2 ,TP6D1 ;
  wire  TP6D0 ,TP5D3 ,TP5D2 ,TP5D1 ,TP5D0 ,TP4D3 ,TP4D2 ,TP4D1 ,TP4D0 ;
  wire  TP3D3 ,TP3D2 ,TP3D1 ,TP3D0 ,TP2D3 ,TP2D2 ,TP2D1 ,TP2D0 ,TP1D3 ;
  wire  TP1D2 ,TP1D1 ,TP1D0 ,CLK30MHZ ,EROMRDB ,EROMCSB ,EROMPA2 ,EROMCLK ,EROMPA17 ;
  wire  EROMPA16 ,EROMPA15 ,EROMPA14 ,EROMPA13 ,EROMPA12 ,EROMPA11 ,EROMPA10 ,EROMPA9 ,EROMPD3 ;
  wire  EROMPA8 ,EROMPD2 ,EROMPA7 ,EROMPD1 ,EROMPA6 ,EROMPD0 ,EROMPA5 ,EROMPA4 ,EROMPA3 ;
  wire  EROMPA1 ,EROMPA0 ,RDCLKP1_OUT ,EXA_OUT ,WWR_OUT ,CER_OUT ,SER_OUT ,EXER_OUT ,MRG00_OUT ;
  wire  MRG01_OUT ,MRG10_OUT ,MRG11_OUT ,MRG12_OUT ,DIS_OUT ,READ_OUT ,FCLK_OUT ,PROGI_OUT ,BFA_OUT ;
  wire  EROMPD31 ,EROMPD23 ,EROMPD15 ,EROMPD30 ,EROMPD22 ,EROMPD14 ,EROMPD29 ,EROMPD28 ,EROMPD27 ;
  wire  EROMPD19 ,EROMPD26 ,EROMPD18 ,EROMPD25 ,EROMPD17 ,EROMPD24 ,EROMPD16 ,EROMPD21 ,EROMPD13 ;
  wire  EROMPD20 ,EROMPD12 ,EROMPD11 ,EROMPD10 ,EROMPD9 ,EROMPD8 ,EROMPD7 ,EROMPD6 ,EROMPD5 ;
  wire  EROMPD4 ,BTFLG ,TMSPMD ,TMBTSEL ,ICETMSPMD ,ICETMBTSEL ,RESB ,USBCLK ,USBRD_B ;
  wire  USBWR0_B ,USBA21 ,USBA20 ,WAITOR ,USBA19 ,USBA4 ,USBA3 ,USBA2 ,USBWAIT_B ;
  wire  USBD15 ,USBD14 ,USBD13 ,USBD12 ,USBD11 ,USBD10 ,USBD9 ,USBD8 ,USBD7 ;
  wire  USBD6 ,USBD5 ,USBD4 ,USBD3 ,USBD2 ,USBD1 ,USBD0 ,ICESYSRES_B ,ICECPURES_B ;
  wire  RESET_B ,EVAOSCMCLK ,EVAOSCRCLK1 ,EVAOSCRCLK2 ,EVAOSCRCLK3 ,TMEMA16 ,TMEMA15 ,TMEMA13 ,TMEMA12 ;
  wire  TMEMA11 ,TMEMA10 ,TMEMA9 ,TMEMD3 ,TMEMA8 ,TMEMD2 ,TMEMA7 ,TMEMD1 ,TMEMA6 ;
  wire  TMEMD0 ,TMEMA5 ,TMEMA4 ,TMEMA3 ,TMEMA2 ,TMEMA1 ,TMEMA0 ,TMEMCS_B ,TMEMRD_B ;
  wire  TMEMWR_B ,TMEMCLK2 ,TMEMCLK1 ,TMEMCLK0 ,TMEMD107 ,TMEMD106 ,TMEMD105 ,TMEMD104 ,TMEMD103 ;
  wire  TMEMD102 ,TMEMD101 ,TMEMD100 ,TMEMD99 ,TMEMD98 ,TMEMD97 ,TMEMD89 ,TMEMD96 ,TMEMD88 ;
  wire  TMEMD95 ,TMEMD87 ,TMEMD79 ,TMEMD94 ,TMEMD86 ,TMEMD78 ,TMEMD93 ,TMEMD85 ,TMEMD77 ;
  wire  TMEMD69 ,TMEMD92 ,TMEMD84 ,TMEMD76 ,TMEMD68 ,TMEMD91 ,TMEMD83 ,TMEMD75 ,TMEMD67 ;
  wire  TMEMD59 ,TMEMD90 ,TMEMD82 ,TMEMD74 ,TMEMD66 ,TMEMD58 ,TMEMD81 ,TMEMD73 ,TMEMD65 ;
  wire  TMEMD57 ,TMEMD49 ,TMEMD80 ,TMEMD72 ,TMEMD64 ,TMEMD56 ,TMEMD48 ,TMEMD71 ,TMEMD63 ;
  wire  TMEMD55 ,TMEMD47 ,TMEMD39 ,TMEMD70 ,TMEMD62 ,TMEMD54 ,TMEMD46 ,TMEMD38 ,TMEMD61 ;
  wire  TMEMD53 ,TMEMD45 ,TMEMD37 ,TMEMD29 ,TMEMD60 ,TMEMD52 ,TMEMD44 ,TMEMD36 ,TMEMD28 ;
  wire  TMEMD51 ,TMEMD43 ,TMEMD35 ,TMEMD27 ,TMEMD19 ,TMEMD50 ,TMEMD42 ,TMEMD34 ,TMEMD26 ;
  wire  TMEMD18 ,TMEMD41 ,TMEMD33 ,TMEMD25 ,TMEMD17 ,TMEMD40 ,TMEMD32 ,TMEMD24 ,TMEMD16 ;
  wire  TMEMD31 ,TMEMD23 ,TMEMD15 ,TMEMD30 ,TMEMD22 ,TMEMD14 ,TMEMD21 ,TMEMD13 ,TMEMD20 ;
  wire  TMEMD12 ,TMEMD11 ,TMEMD10 ,TMEMD9 ,TMEMD8 ,TMEMD7 ,TMEMD6 ,TMEMD5 ,TMEMD4 ;
  wire  TCCONNECT_B ,EACONNECT_B ,TVDDON ,TVDDSEL ,LEDTVDD_B ,LEDCLOCK_B ,LEDRUN_B ,LEDRESET_B ,LEDSTANDBY_B ;
  wire  LEDWAIT_B ,DCE0 ,DCLKSEL1 ,DCER ,DSER ,DWWR ,DWED ,DMRG00 ,DMRG01 ;
  wire  DMRG10 ,DMRG11 ,DMRG12 ,DREAD ,FLMA4 ,AF19 ,AF18 ,AF17 ,DA13 ;
  wire  AF16 ,DA12 ,AF15 ,DA11 ,AF14 ,DA10 ,AF13 ,AF12 ,AF11 ;
  wire  AF10 ,AF9 ,DA7 ,AF8 ,DA6 ,AF5 ,DA3 ,AF4 ,DA2 ;
  wire  AF3 ,DA1 ,AF2 ,DA0 ,AF1 ,AF0 ,DRDCLK ,DRDCLKC1 ,DA9 ;
  wire  DA8 ,DRO11 ,DRO10 ,DRO9 ,DRO8 ,DRO7 ,DRO6 ,DRO5 ,DRO4 ;
  wire  DRO3 ,DRO2 ,DRO1 ,DRO0 ,DDIS_OUT ,ICEDOT26 ,ICEDOT18 ,ICEDOU30 ,ICEDOU22 ;
  wire  ICEDOU14 ,DRDCLKP1_OUT ,DWWR_OUT ,DCER_OUT ,DSER_OUT ,DMRG00_OUT ,DMRG01_OUT ,DMRG10_OUT ,DMRG11_OUT ;
  wire  DMRG12_OUT ,DREAD_OUT ,DFCLK_OUT ,SLDFLASH ,LOCK240FAIL ,CLK240M ,CLK120M ,BFBRKSEL ,ICEFLERRC ;
  wire  EICESYSRES_B ,ICEIFA_PRE31 ,ICEIFA_PRE23 ,ICEIFA_PRE15 ,ICEIFA_PRE30 ,ICEIFA_PRE22 ,ICEIFA_PRE14 ,ICEIFA_PRE29 ,ICEIFA_PRE28 ;
  wire  ICEIFA_PRE27 ,ICEIFA_PRE19 ,ICEIFA_PRE26 ,ICEIFA_PRE18 ,ICEIFA_PRE25 ,ICEIFA_PRE17 ,ICEIFA_PRE24 ,ICEIFA_PRE16 ,ICEIFA_PRE21 ;
  wire  ICEIFA_PRE13 ,ICEIFA_PRE20 ,ICEIFA_PRE12 ,ICEIFA_PRE11 ,ICEIFA_PRE10 ,ICEIFA_PRE9 ,ICEIFA_PRE8 ,ICEIFA_PRE7 ,ICEIFA_PRE6 ;
  wire  ICEIFA_PRE5 ,ICEIFA_PRE4 ,ICEIFA_PRE3 ,ICEIFA_PRE2 ,ICEDI_PRE0 ,ICEWR_PRE ,EICECPURES_B ,BRKFAIL14 ,BRKTMOVR ;
  wire  BRKTMOVC0 ,BRKTMOVC1 ,BRKTMOVN0 ,BRKTMOVN1 ,BRKSNAP2 ,BRKSNAP1 ,BRKSNAP0 ,BRKEDMM3 ,BRKEDMM2 ;
  wire  BRKEDMM1 ,BRKEDMM0 ,ETCCONNECT_B ,EEACONNECT_B ,ETVDDSEL ,ELEDTVDD_B ,ELEDCLOCK_B ,ELEDRUN_B ,ELEDRESET_B ;
  wire  ELEDSTANDBY_B ,ELEDWAIT_B ,SWAP ,ADDRICE0 ,UP ,ADDRICE1 ,ADDRICE2 ,ADDRICE3 ,ADDRICE4 ;
  wire  ADDRICE5 ,ADDRICE6 ,ADDRICE7 ,ADDRICE8 ,ADDRICE9 ,ADDRICE10 ,ADDRICE11 ,TVDDSELB ,ICEDOE31 ;
  wire  ICEDOE23 ,ICEDOE15 ,ICEDOD27 ,ICEDOD19 ,ICEDOF11 ,ICEDOE30 ,ICEDOE22 ,ICEDOE14 ,ICEDOD26 ;
  wire  ICEDOD18 ,ICEDOF10 ,ICEDOE29 ,ICEDOF25 ,ICEDOF17 ,ICEDOG21 ,ICEDOG13 ,ICEDOE28 ,ICEDOF24 ;
  wire  ICEDOF16 ,ICEDOG20 ,ICEDOG12 ,ICEDOE27 ,ICEDOE19 ,ICEDOF31 ,ICEDOF23 ,ICEDOF15 ,ICEDOG11 ;
  wire  ICEDOE26 ,ICEDOE18 ,ICEDOF30 ,ICEDOF22 ,ICEDOF14 ,ICEDOG10 ,ICEDOE25 ,ICEDOE17 ,ICEDOD29 ;
  wire  ICEDOF21 ,ICEDOF13 ,ICEDOE24 ,ICEDOE16 ,ICEDOD28 ,ICEDOF20 ,ICEDOF12 ,ICEDOE9 ,ICEDOF7 ;
  wire  ICEDOG5 ,ICEDOH3 ,ICEDOE8 ,ICEDOF6 ,ICEDOG4 ,ICEDOH2 ,ICEDOE7 ,ICEDOD9 ,ICEDOF5 ;
  wire  ICEDOG3 ,ICEDOH1 ,ICEDOE6 ,ICEDOD8 ,ICEDOF4 ,ICEDOG2 ,ICEDOH0 ,HOSTIFMDR15 ,HOSTIFMDR14 ;
  wire  HOSTIFMDR13 ,HOSTIFMDR12 ,HOSTIFMDR11 ,HOSTIFMDR10 ,HOSTIFMDR9 ,HOSTIFMDR8 ,HOSTIFMDR7 ,HOSTIFMDR6 ,HOSTIFMDR5 ;
  wire  HOSTIFMDR4 ,HOSTIFMDR3 ,HOSTIFMDR2 ,HOSTIFMDR1 ,HOSTIFMDR0 ,ICEDOF29 ,ICEDOG25 ,ICEDOG17 ,ICEDOH21 ;
  wire  ICEDOH13 ,ICEDOF28 ,ICEDOG24 ,ICEDOG16 ,ICEDOH20 ,ICEDOH12 ,ICEDOF27 ,ICEDOF19 ,ICEDOG31 ;
  wire  ICEDOG23 ,ICEDOG15 ,ICEDOH11 ,ICEDOF26 ,ICEDOF18 ,ICEDOG30 ,ICEDOG22 ,ICEDOG14 ,ICEDOH10 ;
  wire  ICEDOF9 ,ICEDOG7 ,ICEDOH5 ,ICEDOJ1 ,ICEDOF8 ,ICEDOG6 ,ICEDOH4 ,ICEDOJ0 ,BRKMDR15 ;
  wire  BRKMDR14 ,BRKMDR13 ,BRKMDR12 ,BRKMDR11 ,BRKMDR10 ,BRKMDR9 ,BRKMDR8 ,BRKMDR7 ,BRKMDR6 ;
  wire  BRKMDR5 ,BRKMDR4 ,BRKMDR3 ,BRKMDR2 ,ICEDOG29 ,ICEDOH25 ,ICEDOH17 ,ICEDOG28 ,ICEDOH24 ;
  wire  ICEDOH16 ,ICEDOG27 ,ICEDOG19 ,ICEDOH31 ,ICEDOH23 ,ICEDOH15 ,ICEDOG26 ,ICEDOG18 ,ICEDOH30 ;
  wire  ICEDOH22 ,ICEDOH14 ,ICEDOG9 ,ICEDOK1 ,ICEDOH7 ,ICEDOJ3 ,ICEDOG8 ,ICEDOK0 ,ICEDOH6 ;
  wire  ICEDOJ2 ,ICEDOK31 ,ICEDOK23 ,ICEDOK15 ,ICEDOJ27 ,ICEDOJ19 ,ICEDOL11 ,ICEDOK30 ,ICEDOK22 ;
  wire  ICEDOK14 ,ICEDOJ26 ,ICEDOJ18 ,ICEDOL10 ,ICEDOK29 ,ICEDOM21 ,ICEDOM13 ,ICEDOL25 ,ICEDOL17 ;
  wire  ICEDOK28 ,ICEDOM20 ,ICEDOM12 ,ICEDOL24 ,ICEDOL16 ,ICEDOK27 ,ICEDOK19 ,ICEDOM11 ,ICEDOL31 ;
  wire  ICEDOL23 ,ICEDOL15 ,ICEDOK26 ,ICEDOK18 ,ICEDOM10 ,ICEDOL30 ,ICEDOL22 ,ICEDOL14 ,ICEDOK25 ;
  wire  ICEDOK17 ,ICEDOJ29 ,ICEDOL21 ,ICEDOL13 ,ICEDOK24 ,ICEDOK16 ,ICEDOJ28 ,ICEDOL20 ,ICEDOL12 ;
  wire  ICEDOK21 ,ICEDOK13 ,ICEDOJ25 ,ICEDOJ17 ,ICEDOK20 ,ICEDOK12 ,ICEDOJ24 ,ICEDOJ16 ,ICEDOK11 ;
  wire  ICEDOJ31 ,ICEDOJ23 ,ICEDOJ15 ,ICEDOK10 ,ICEDOJ30 ,ICEDOJ22 ,ICEDOJ14 ,ICEDOK9 ,ICEDON3 ;
  wire  ICEDOM5 ,ICEDOL7 ,ICEDOK8 ,ICEDON2 ,ICEDOM4 ,ICEDOL6 ,ICEDOK7 ,ICEDOJ9 ,ICEDON1 ;
  wire  ICEDOM3 ,ICEDOL5 ,ICEDOK6 ,ICEDOJ8 ,ICEDON0 ,ICEDOM2 ,ICEDOL4 ,ICEDOK5 ,ICEDOJ7 ;
  wire  ICEDOM1 ,ICEDOL3 ,ICEDOK4 ,ICEDOJ6 ,ICEDOM0 ,ICEDOL2 ,ICEDOK3 ,ICEDOH9 ,ICEDOJ5 ;
  wire  ICEDOL1 ,ICEDOK2 ,ICEDOH8 ,ICEDOJ4 ,ICEDOL0 ,ICEDOH29 ,ICEDOJ21 ,ICEDOJ13 ,ICEDOH28 ;
  wire  ICEDOJ20 ,ICEDOJ12 ,ICEDOH27 ,ICEDOH19 ,ICEDOJ11 ,ICEDOH26 ,ICEDOH18 ,ICEDOJ10 ,ICEDOQ29 ;
  wire  ICEDOS21 ,ICEDOS13 ,ICEDOR25 ,ICEDOR17 ,ICEDOQ28 ,ICEDOS20 ,ICEDOS12 ,ICEDOR24 ,ICEDOR16 ;
  wire  ICEDOQ27 ,ICEDOQ19 ,ICEDOS11 ,ICEDOR31 ,ICEDOR23 ,ICEDOR15 ,ICEDOQ26 ,ICEDOQ18 ,ICEDOS10 ;
  wire  ICEDOR30 ,ICEDOR22 ,ICEDOR14 ,ICEDOQ9 ,ICEDOS5 ,ICEDOT3 ,ICEDOR7 ,ICEDOU1 ,ICEDOQ8 ;
  wire  ICEDOS4 ,ICEDOT2 ,ICEDOR6 ,ICEDOU0 ,ICEDON31 ,ICEDON23 ,ICEDON15 ,ICEDOM27 ,ICEDOM19 ;
  wire  ICEDON30 ,ICEDON22 ,ICEDON14 ,ICEDOM26 ,ICEDOM18 ,ICEDON25 ,ICEDON17 ,ICEDOM29 ,ICEDON24 ;
  wire  ICEDON16 ,ICEDOM28 ,ICEDON21 ,ICEDON13 ,ICEDOM25 ,ICEDOM17 ,ICEDOL29 ,ICEDON20 ,ICEDON12 ;
  wire  ICEDOM24 ,ICEDOM16 ,ICEDOL28 ,ICEDON11 ,ICEDOM31 ,ICEDOM23 ,ICEDOM15 ,ICEDOL27 ,ICEDOL19 ;
  wire  ICEDON10 ,ICEDOM30 ,ICEDOM22 ,ICEDOM14 ,ICEDOL26 ,ICEDOL18 ,ICEDOS31 ,ICEDOS23 ,ICEDOS15 ;
  wire  ICEDOT11 ,ICEDOR27 ,ICEDOR19 ,ICEDOS30 ,ICEDOS22 ,ICEDOS14 ,ICEDOT10 ,ICEDOR26 ,ICEDOR18 ;
  wire  ICEDOS29 ,ICEDOT25 ,ICEDOT17 ,ICEDOU21 ,ICEDOU13 ,ICEDOS28 ,ICEDOT24 ,ICEDOT16 ,ICEDOU20 ;
  wire  ICEDOU12 ,ICEDOS27 ,ICEDOS19 ,ICEDOT31 ,ICEDOT23 ,ICEDOT15 ,ICEDOU11 ,ICEDOS26 ,ICEDOS18 ;
  wire  ICEDOT30 ,ICEDOT22 ,ICEDOT14 ,ICEDOU10 ,ICEDOS25 ,ICEDOS17 ,ICEDOT21 ,ICEDOT13 ,ICEDOR29 ;
  wire  ICEDOS24 ,ICEDOS16 ,ICEDOT20 ,ICEDOT12 ,ICEDOR28 ,ICEDOS9 ,ICEDOT7 ,ICEDOU5 ,ICEDOS8 ;
  wire  ICEDOT6 ,ICEDOU4 ,ICEDOS7 ,ICEDOT5 ,ICEDOR9 ,ICEDOU3 ,ICEDOS6 ,ICEDOT4 ,ICEDOR8 ;
  wire  ICEDOU2 ,ICEDOT29 ,ICEDOU25 ,ICEDOU17 ,ICEDOT28 ,ICEDOU24 ,ICEDOU16 ,ICEDOT27 ,ICEDOT19 ;
  wire  ICEDOU31 ,ICEDOU23 ,ICEDOU15 ,ICEDOT9 ,ICEDOU7 ,ICEDOT8 ,ICEDOU6 ,TI0D3 ,TI0D2 ;
  wire  TI0D1 ,TAG29 ,TI0D0 ,TAG28 ,TI1D3 ,TI1D2 ,TI1D1 ,TI2D3 ,TI2D2 ;
  wire  TI2D1 ,TI2D0 ,TI4D3 ,TI4D2 ,TI4D1 ,TI5D3 ,TI5D2 ,TI5D1 ,TI5D0 ;
  wire  TI6D3 ,TI6D2 ,TI6D1 ,TI6D0 ,TI7D3 ,TI7D2 ,TI7D1 ,TI7D0 ,TI8D3 ;
  wire  TI8D2 ,TI8D1 ,TI8D0 ,TI9D3 ,TI9D2 ,TI9D1 ,TI9D0 ,TI10D3 ,TI10D2 ;
  wire  TI10D1 ,TI10D0 ,TI11D3 ,TI11D2 ,TI11D1 ,TI11D0 ,MONITRC ,TAG31 ,TAG23 ;
  wire  TAG15 ,TAG30 ,TAG22 ,TAG14 ,TAG27 ,TAG19 ,TAG26 ,TAG18 ,TAG25 ;
  wire  TAG17 ,TAG24 ,TAG16 ,TAG9 ,TAG7 ,TAG6 ,TAGOVF ,EVD14 ,FLMA0 ;
  wire  EVD06 ,EVD13 ,EVD05 ,EVD12 ,ICERD ,EVD04 ,EVD11 ,EVD03 ,BRKTMOT0 ;
  wire  BRKTMOT1 ,EROMWAIT ,MEMMDR15 ,MEMMDR14 ,MEMMDR13 ,MEMMDR12 ,MEMMDR11 ,MEMMDR10 ,MEMMDR9 ;
  wire  MEMMDR8 ,MEMMDR7 ,MEMMDR5 ,MEMMDR4 ,MEMMDR3 ,MEMMDR2 ,MEMMDR1 ,MEMMDR0 ,FLMA15 ;
  wire  FLMA14 ,FLMA13 ,FLMA12 ,FLMA11 ,FLMA10 ,FLMA9 ,FLMA8 ,FLMA7 ,FLMA5 ;
  wire  FLMA3 ,EVD09 ,FLMA2 ,EVD08 ,FLMA1 ,EVD07 ,MAAOUT ,SELFMODE ,SELFMODEDBG ;
  wire  FAILMK12 ,BRKFAIL12 ,BFBRKPID31 ,BFBRKPID23 ,BFBRKPID15 ,BFBRKPID30 ,BFBRKPID22 ,BFBRKPID14 ,BFBRKPID29 ;
  wire  BFBRKPID28 ,BFBRKPID27 ,BFBRKPID19 ,BFBRKPID26 ,BFBRKPID18 ,BFBRKPID25 ,BFBRKPID17 ,BFBRKPID24 ,BFBRKPID16 ;
  wire  BFBRKPID21 ,BFBRKPID13 ,BFBRKPID20 ,BFBRKPID12 ,BFBRKPID11 ,BFBRKPID10 ,BFBRKPID9 ,BFBRKPID8 ,BFBRKPID7 ;
  wire  BFBRKPID6 ,BFBRKPID5 ,BFBRKPID4 ,BFBRKPID3 ,BFBRKPID2 ,BFBRKPID1 ,BFBRKPID0 ,ICEDOU29 ,ICEDOU28 ;
  wire  ICEDOU27 ,ICEDOU19 ,ICEDOU26 ,ICEDOU18 ,ICEDOU9 ,ICEDOU8 ,ICEIFA_PRE1 ,ICEIFA_PRE0 ,ICEDI_PRE31 ;
  wire  ICEDI_PRE23 ,ICEDI_PRE15 ,ICEDI_PRE30 ,ICEDI_PRE22 ,ICEDI_PRE14 ,ICEDI_PRE29 ,ICEDI_PRE28 ,ICEDI_PRE27 ,ICEDI_PRE19 ;
  wire  ICEDI_PRE26 ,ICEDI_PRE18 ,ICEDI_PRE25 ,ICEDI_PRE17 ,ICEDI_PRE24 ,ICEDI_PRE16 ,ICEDI_PRE21 ,ICEDI_PRE13 ,ICEDI_PRE20 ;
  wire  ICEDI_PRE12 ,ICEDI_PRE11 ,ICEDI_PRE10 ,ICEDI_PRE9 ,ICEDI_PRE8 ,ICEDI_PRE7 ,ICEDI_PRE6 ,ICEDI_PRE5 ,ICEDI_PRE4 ;
  wire  ICEDI_PRE3 ,ICEDI_PRE2 ,ICEDI_PRE1 ,ICERD_PRE ,SVMODUSER ,PSEUDORES ,TRACEMDR1 ,ICEMSKPOC ,ICEMSKTRST ;
  wire  ICEMSKICE ,ICEMSKTRSTFLG ,ICERESB ,TARRESB_NORM ,BRKFAIL0 ,BRKFAIL1 ,BRKFAIL2 ,BRKFAIL3 ,BRKFAIL4 ;
  wire  BRKFAIL5 ,BRKFAIL6 ,BRKFAIL7 ,BRKFAIL8 ,BRKFAIL9 ,BRKFAIL10 ,BRKFAIL11 ,BRKFAIL13 ,BRKFAIL15 ;
  wire  BRKEVTF0 ,BRKEVTF1 ,BRKEVTF2 ,BRKEVTF3 ,BRKEVTF4 ,BRKEVTF5 ,BRKEVTF6 ,BRKEVTF7 ,BRKEVTA0 ;
  wire  BRKEVTA1 ,BRKEVTA2 ,BRKEVTA3 ,BRKEVTA4 ,BRKEVTA5 ,BRKEVTA6 ,BRKEVTA7 ,BRKEVTL0 ,BRKEVTL1 ;
  wire  BRKTRAFL ,BRKTRADY ,STEP ,TRACEMDR15 ,TRACEMDR14 ,TRACEMDR13 ,TRACEMDR12 ,TRACEMDR11 ,TRACEMDR10 ;
  wire  TRACEMDR9 ,TRACEMDR8 ,TRACEMDR7 ,TRACEMDR6 ,TRACEMDR5 ,TRACEMDR4 ,TRACEMDR3 ,TRACEMDR2 ,TRACEMDR0 ;
  wire  SELEXMPC ,SELRAMPC ,SELROMPC ,SELBRAMPC ,SELBFAPC ,EVD01 ,EVD02 ,EVD10 ,TRCON ;
  wire  TRCMD ,TMEMWAIT ,EXMAPOUT ,STATEMDR15 ,STATEMDR14 ,STATEMDR13 ,STATEMDR12 ,STATEMDR11 ,STATEMDR10 ;
  wire  STATEMDR9 ,STATEMDR8 ,STATEMDR7 ,STATEMDR6 ,STATEMDR5 ,STATEMDR4 ,STATEMDR3 ,STATEMDR2 ,STATEMDR1 ;
  wire  STATEMDR0 ,DFMDR15 ,DFMDR14 ,DFMDR13 ,DFMDR12 ,DFMDR11 ,DFMDR10 ,DFMDR9 ,DFMDR8 ;
  wire  DFMDR7 ,DFMDR6 ,DFMDR5 ,DFMDR4 ,DFMDR3 ,DFMDR2 ,DFMDR0 ,ICEFLERRD ;


  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/iirl78timetagv1.v
  IIRL78TIMETAGV1 timetagv2 (
   .ICEIFA31 ( ICEIFA31 ) ,.ICEIFA23 ( ICEIFA23 ) ,.ICEIFA15 ( ICEIFA15 ) ,.ICEIFA30 ( ICEIFA30 ) ,.ICEIFA22 ( ICEIFA22 ) ,.ICEIFA14 ( ICEIFA14 ) ,.ICEIFA29 ( ICEIFA29 )
 ,.ICEIFA28 ( ICEIFA28 ) ,.ICEIFA27 ( ICEIFA27 ) ,.ICEIFA19 ( ICEIFA19 ) ,.ICEIFA26 ( ICEIFA26 ) ,.ICEIFA18 ( ICEIFA18 ) ,.ICEIFA25 ( ICEIFA25 )
 ,.ICEIFA17 ( ICEIFA17 ) ,.ICEIFA24 ( ICEIFA24 ) ,.ICEIFA16 ( ICEIFA16 ) ,.ICEIFA21 ( ICEIFA21 ) ,.ICEIFA13 ( ICEIFA13 ) ,.ICEIFA20 ( ICEIFA20 )
 ,.ICEIFA12 ( ICEIFA12 ) ,.ICEIFA11 ( ICEIFA11 ) ,.ICEIFA10 ( ICEIFA10 ) ,.ICEIFA9 ( ICEIFA9 ) ,.ICEIFA8 ( ICEIFA8 ) ,.ICEIFA7 ( ICEIFA7 )
 ,.ICEIFA6 ( ICEIFA6 ) ,.ICEIFA5 ( ICEIFA5 ) ,.ICEIFA4 ( ICEIFA4 ) ,.ICEIFA3 ( ICEIFA3 ) ,.ICEIFA2 ( ICEIFA2 ) ,.ICEIFA1 ( ICEIFA1 )
 ,.ICEIFA0 ( ICEIFA0 ) ,.ICEDI31 ( ICEDI31 ) ,.ICEDI23 ( ICEDI23 ) ,.ICEDI15 ( ICEDI15 ) ,.ICEDI30 ( ICEDI30 ) ,.ICEDI22 ( ICEDI22 )
 ,.ICEDI14 ( ICEDI14 ) ,.ICEDI29 ( ICEDI29 ) ,.ICEDI28 ( ICEDI28 ) ,.ICEDI27 ( ICEDI27 ) ,.ICEDI19 ( ICEDI19 ) ,.ICEDI26 ( ICEDI26 )
 ,.ICEDI18 ( ICEDI18 ) ,.ICEDI25 ( ICEDI25 ) ,.ICEDI17 ( ICEDI17 ) ,.ICEDI24 ( ICEDI24 ) ,.ICEDI16 ( ICEDI16 ) ,.ICEDI21 ( ICEDI21 )
 ,.ICEDI13 ( ICEDI13 ) ,.ICEDI20 ( ICEDI20 ) ,.ICEDI12 ( ICEDI12 ) ,.ICEDI11 ( ICEDI11 ) ,.ICEDI10 ( ICEDI10 ) ,.ICEDI9 ( ICEDI9 )
 ,.ICEDI8 ( ICEDI8 ) ,.ICEDI7 ( ICEDI7 ) ,.ICEDI6 ( ICEDI6 ) ,.ICEDI5 ( ICEDI5 ) ,.ICEDI4 ( ICEDI4 ) ,.ICEDI3 ( ICEDI3 )
 ,.ICEDI2 ( ICEDI2 ) ,.ICEDI1 ( ICEDI1 ) ,.ICEDI0 ( ICEDI0 ) ,.ICEWR ( ICEWR ) ,.ICEDOR31 ( ICEDOR31 ) ,.ICEDOR23 ( ICEDOR23 )
 ,.ICEDOR15 ( ICEDOR15 ) ,.ICEDOR30 ( ICEDOR30 ) ,.ICEDOR22 ( ICEDOR22 ) ,.ICEDOR14 ( ICEDOR14 ) ,.ICEDOR29 ( ICEDOR29 ) ,.ICEDOR28 ( ICEDOR28 )
 ,.ICEDOR27 ( ICEDOR27 ) ,.ICEDOR19 ( ICEDOR19 ) ,.ICEDOR26 ( ICEDOR26 ) ,.ICEDOR18 ( ICEDOR18 ) ,.ICEDOR25 ( ICEDOR25 ) ,.ICEDOR17 ( ICEDOR17 )
 ,.ICEDOR24 ( ICEDOR24 ) ,.ICEDOR16 ( ICEDOR16 ) ,.ICEDOR21 ( ICEDOR21 ) ,.ICEDOR13 ( ICEDOR13 ) ,.ICEDOR20 ( ICEDOR20 ) ,.ICEDOR12 ( ICEDOR12 )
 ,.ICEDOR11 ( ICEDOR11 ) ,.ICEDOR10 ( ICEDOR10 ) ,.ICEDOR9 ( ICEDOR9 ) ,.ICEDOR8 ( ICEDOR8 ) ,.ICEDOR7 ( ICEDOR7 ) ,.ICEDOR6 ( ICEDOR6 )
 ,.ICEDOR5 ( ICEDOR5 ) ,.ICEDOR4 ( ICEDOR4 ) ,.ICEDOR3 ( ICEDOR3 ) ,.ICEDOR2 ( ICEDOR2 ) ,.ICEDOR1 ( ICEDOR1 ) ,.ICEDOR0 ( ICEDOR0 )
 ,.BASECK ( BASECK ) ,.SYSRSOUTB ( SYSRSOUTB ) ,.SVMODI ( SVMODI ) ,.MONITRC ( MONITRC ) ,.TAG31 ( TAG31 ) ,.TAG23 ( TAG23 )
 ,.TAG15 ( TAG15 ) ,.TAG30 ( TAG30 ) ,.TAG22 ( TAG22 ) ,.TAG14 ( TAG14 ) ,.TAG29 ( TAG29 ) ,.TAG28 ( TAG28 )
 ,.TAG27 ( TAG27 ) ,.TAG19 ( TAG19 ) ,.TAG26 ( TAG26 ) ,.TAG18 ( TAG18 ) ,.TAG25 ( TAG25 ) ,.TAG17 ( TAG17 )
 ,.TAG24 ( TAG24 ) ,.TAG16 ( TAG16 ) ,.TAG21 ( TAG21 ) ,.TAG13 ( TAG13 ) ,.TAG20 ( TAG20 ) ,.TAG12 ( TAG12 )
 ,.TAG11 ( TAG11 ) ,.TAG10 ( TAG10 ) ,.TAG9 ( TAG9 ) ,.TAG8 ( TAG8 ) ,.TAG7 ( TAG7 ) ,.TAG6 ( TAG6 )
 ,.TAG5 ( TAG5 ) ,.TAG4 ( TAG4 ) ,.TAG3 ( TAG3 ) ,.TAG2 ( TAG2 ) ,.TAG1 ( TAG1 ) ,.TAG0 ( TAG0 )
 ,.TAGOVF ( TAGOVF ) ,.CLK240M ( CLK240M )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/iirl78timerv1.v
  IIRL78TIMERV1 timerv2 (
   .ICEDO31 ( ICEDON31 ) ,.ICEDO23 ( ICEDON23 ) ,.ICEDO15 ( ICEDON15 ) ,.ICEDO30 ( ICEDON30 ) ,.ICEDO22 ( ICEDON22 ) ,.ICEDO14 ( ICEDON14 ) ,.ICEDO29 ( ICEDON29 )
 ,.ICEDO28 ( ICEDON28 ) ,.ICEDO27 ( ICEDON27 ) ,.ICEDO19 ( ICEDON19 ) ,.ICEDO26 ( ICEDON26 ) ,.ICEDO18 ( ICEDON18 ) ,.ICEDO25 ( ICEDON25 )
 ,.ICEDO17 ( ICEDON17 ) ,.ICEDO24 ( ICEDON24 ) ,.ICEDO16 ( ICEDON16 ) ,.ICEDO21 ( ICEDON21 ) ,.ICEDO13 ( ICEDON13 ) ,.ICEDO20 ( ICEDON20 )
 ,.ICEDO12 ( ICEDON12 ) ,.ICEDO11 ( ICEDON11 ) ,.ICEDO10 ( ICEDON10 ) ,.ICEDO9 ( ICEDON9 ) ,.ICEDO8 ( ICEDON8 ) ,.ICEDO7 ( ICEDON7 )
 ,.ICEDO6 ( ICEDON6 ) ,.ICEDO5 ( ICEDON5 ) ,.ICEDO4 ( ICEDON4 ) ,.ICEDO3 ( ICEDON3 ) ,.ICEDO2 ( ICEDON2 ) ,.ICEDO1 ( ICEDON1 )
 ,.ICEDO0 ( ICEDON0 ) ,.ICEIFA31 ( ICEIFA31 ) ,.ICEIFA23 ( ICEIFA23 ) ,.ICEIFA15 ( ICEIFA15 ) ,.ICEIFA30 ( ICEIFA30 ) ,.ICEIFA22 ( ICEIFA22 )
 ,.ICEIFA14 ( ICEIFA14 ) ,.ICEIFA29 ( ICEIFA29 ) ,.ICEIFA28 ( ICEIFA28 ) ,.ICEIFA27 ( ICEIFA27 ) ,.ICEIFA19 ( ICEIFA19 ) ,.ICEIFA26 ( ICEIFA26 )
 ,.ICEIFA18 ( ICEIFA18 ) ,.ICEIFA25 ( ICEIFA25 ) ,.ICEIFA17 ( ICEIFA17 ) ,.ICEIFA24 ( ICEIFA24 ) ,.ICEIFA16 ( ICEIFA16 ) ,.ICEIFA21 ( ICEIFA21 )
 ,.ICEIFA13 ( ICEIFA13 ) ,.ICEIFA20 ( ICEIFA20 ) ,.ICEIFA12 ( ICEIFA12 ) ,.ICEIFA11 ( ICEIFA11 ) ,.ICEIFA10 ( ICEIFA10 ) ,.ICEIFA9 ( ICEIFA9 )
 ,.ICEIFA8 ( ICEIFA8 ) ,.ICEIFA7 ( ICEIFA7 ) ,.ICEIFA6 ( ICEIFA6 ) ,.ICEIFA5 ( ICEIFA5 ) ,.ICEIFA4 ( ICEIFA4 ) ,.ICEIFA3 ( ICEIFA3 )
 ,.ICEIFA2 ( ICEIFA2 ) ,.ICEIFA1 ( ICEIFA1 ) ,.ICEIFA0 ( ICEIFA0 ) ,.ICEDI31 ( ICEDI31 ) ,.ICEDI23 ( ICEDI23 ) ,.ICEDI15 ( ICEDI15 )
 ,.ICEDI30 ( ICEDI30 ) ,.ICEDI22 ( ICEDI22 ) ,.ICEDI14 ( ICEDI14 ) ,.ICEDI29 ( ICEDI29 ) ,.ICEDI28 ( ICEDI28 ) ,.ICEDI27 ( ICEDI27 )
 ,.ICEDI19 ( ICEDI19 ) ,.ICEDI26 ( ICEDI26 ) ,.ICEDI18 ( ICEDI18 ) ,.ICEDI25 ( ICEDI25 ) ,.ICEDI17 ( ICEDI17 ) ,.ICEDI24 ( ICEDI24 )
 ,.ICEDI16 ( ICEDI16 ) ,.ICEDI21 ( ICEDI21 ) ,.ICEDI13 ( ICEDI13 ) ,.ICEDI20 ( ICEDI20 ) ,.ICEDI12 ( ICEDI12 ) ,.ICEDI11 ( ICEDI11 )
 ,.ICEDI10 ( ICEDI10 ) ,.ICEDI9 ( ICEDI9 ) ,.ICEDI8 ( ICEDI8 ) ,.ICEDI7 ( ICEDI7 ) ,.ICEDI6 ( ICEDI6 ) ,.ICEDI5 ( ICEDI5 )
 ,.ICEDI4 ( ICEDI4 ) ,.ICEDI3 ( ICEDI3 ) ,.ICEDI2 ( ICEDI2 ) ,.ICEDI1 ( ICEDI1 ) ,.ICEDI0 ( ICEDI0 ) ,.ICEWR ( ICEWR )
 ,.EVD14 ( EVD14 ) ,.EVD13 ( EVD13 ) ,.EVD12 ( EVD12 ) ,.EVD11 ( EVD11 ) ,.BRKTMOVR ( BRKTMOVR ) ,.BRKTMOVC0 ( BRKTMOVC0 )
 ,.BRKTMOVN0 ( BRKTMOVN0 ) ,.BRKTMOVC1 ( BRKTMOVC1 ) ,.BRKTMOVN1 ( BRKTMOVN1 ) ,.BRKTMOT0 ( BRKTMOT0 ) ,.BRKTMOT1 ( BRKTMOT1 ) ,.BASECK ( BASECK )
 ,.SYSRSOUTB ( SYSRSOUTB ) ,.SVMODI ( SVMODI ) ,.CLK120M ( CLK120M )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/emem-SS3rd.v
  EVA_EMEM emem (
   .WAITMEM ( ICEWAITMEM ) ,.BFBRKCTL ( BFBRKSEL ) ,.CPURESETB ( CPURSOUTB ) ,.CK60MHZ ( CLK60MHZ ) ,.ICEFLERR ( ICEFLERRC ) ,.ICEDO31 ( ICEDOE31 ) ,.ICEDO23 ( ICEDOE23 )
 ,.ICEDO15 ( ICEDOE15 ) ,.ICEDO30 ( ICEDOE30 ) ,.ICEDO22 ( ICEDOE22 ) ,.ICEDO14 ( ICEDOE14 ) ,.ICEDO29 ( ICEDOE29 ) ,.ICEDO28 ( ICEDOE28 )
 ,.ICEDO27 ( ICEDOE27 ) ,.ICEDO19 ( ICEDOE19 ) ,.ICEDO26 ( ICEDOE26 ) ,.ICEDO18 ( ICEDOE18 ) ,.ICEDO25 ( ICEDOE25 ) ,.ICEDO17 ( ICEDOE17 )
 ,.ICEDO24 ( ICEDOE24 ) ,.ICEDO16 ( ICEDOE16 ) ,.ICEDO21 ( ICEDOE21 ) ,.ICEDO13 ( ICEDOE13 ) ,.ICEDO20 ( ICEDOE20 ) ,.ICEDO12 ( ICEDOE12 )
 ,.ICEDO11 ( ICEDOE11 ) ,.ICEDO10 ( ICEDOE10 ) ,.ICEDO9 ( ICEDOE9 ) ,.ICEDO8 ( ICEDOE8 ) ,.ICEDO7 ( ICEDOE7 ) ,.ICEDO6 ( ICEDOE6 )
 ,.ICEDO5 ( ICEDOE5 ) ,.ICEDO4 ( ICEDOE4 ) ,.ICEDO3 ( ICEDOE3 ) ,.ICEDO2 ( ICEDOE2 ) ,.ICEDO1 ( ICEDOE1 ) ,.ICEDO0 ( ICEDOE0 )
 ,.EROMRDB ( EROMRDB ) ,.EROMWRB ( EROMWRB ) ,.EROMCSB ( EROMCSB ) ,.EROMPA2 ( EROMPA2 ) ,.EROMCLK ( EROMCLK ) ,.EROMPA17 ( EROMPA17 )
 ,.EROMPA16 ( EROMPA16 ) ,.EROMPA15 ( EROMPA15 ) ,.EROMPA14 ( EROMPA14 ) ,.EROMPA13 ( EROMPA13 ) ,.EROMPA12 ( EROMPA12 ) ,.EROMPA11 ( EROMPA11 )
 ,.EROMPA10 ( EROMPA10 ) ,.EROMPA9 ( EROMPA9 ) ,.EROMPD3 ( EROMPD3 ) ,.EROMPA8 ( EROMPA8 ) ,.EROMPD2 ( EROMPD2 ) ,.EROMPA7 ( EROMPA7 )
 ,.EROMPD1 ( EROMPD1 ) ,.EROMPA6 ( EROMPA6 ) ,.EROMPD0 ( EROMPD0 ) ,.EROMPA5 ( EROMPA5 ) ,.EROMPA4 ( EROMPA4 ) ,.EROMPA3 ( EROMPA3 )
 ,.EROMPA1 ( EROMPA1 ) ,.EROMPA0 ( EROMPA0 ) ,.EROMPD31 ( EROMPD31 ) ,.EROMPD23 ( EROMPD23 ) ,.EROMPD15 ( EROMPD15 ) ,.EROMPD30 ( EROMPD30 )
 ,.EROMPD22 ( EROMPD22 ) ,.EROMPD14 ( EROMPD14 ) ,.EROMPD29 ( EROMPD29 ) ,.EROMPD28 ( EROMPD28 ) ,.EROMPD27 ( EROMPD27 ) ,.EROMPD19 ( EROMPD19 )
 ,.EROMPD26 ( EROMPD26 ) ,.EROMPD18 ( EROMPD18 ) ,.EROMPD25 ( EROMPD25 ) ,.EROMPD17 ( EROMPD17 ) ,.EROMPD24 ( EROMPD24 ) ,.EROMPD16 ( EROMPD16 )
 ,.EROMPD21 ( EROMPD21 ) ,.EROMPD13 ( EROMPD13 ) ,.EROMPD20 ( EROMPD20 ) ,.EROMPD12 ( EROMPD12 ) ,.EROMPD11 ( EROMPD11 ) ,.EROMPD10 ( EROMPD10 )
 ,.EROMPD9 ( EROMPD9 ) ,.EROMPD8 ( EROMPD8 ) ,.EROMPD7 ( EROMPD7 ) ,.EROMPD6 ( EROMPD6 ) ,.EROMPD5 ( EROMPD5 ) ,.EROMPD4 ( EROMPD4 )
 ,.RDCLKP1_OUT ( RDCLKP1_OUT ) ,.EXA_OUT ( EXA_OUT ) ,.WWR_OUT ( WWR_OUT ) ,.CER_OUT ( CER_OUT ) ,.SER_OUT ( SER_OUT ) ,.EXER_OUT ( EXER_OUT )
 ,.MRG00_OUT ( MRG00_OUT ) ,.MRG01_OUT ( MRG01_OUT ) ,.MRG10_OUT ( MRG10_OUT ) ,.MRG11_OUT ( MRG11_OUT ) ,.MRG12_OUT ( MRG12_OUT ) ,.DIS_OUT ( DIS_OUT )
 ,.READ_OUT ( READ_OUT ) ,.FCLK_OUT ( FCLK_OUT ) ,.PROGI_OUT ( PROGI_OUT ) ,.BFA_OUT ( BFA_OUT ) ,.ICEIFA31 ( ICEIFA31 ) ,.ICEIFA23 ( ICEIFA23 )
 ,.ICEIFA15 ( ICEIFA15 ) ,.ICEIFA30 ( ICEIFA30 ) ,.ICEIFA22 ( ICEIFA22 ) ,.ICEIFA14 ( ICEIFA14 ) ,.ICEIFA29 ( ICEIFA29 ) ,.ICEIFA28 ( ICEIFA28 )
 ,.ICEIFA27 ( ICEIFA27 ) ,.ICEIFA19 ( ICEIFA19 ) ,.ICEIFA26 ( ICEIFA26 ) ,.ICEIFA18 ( ICEIFA18 ) ,.ICEIFA25 ( ICEIFA25 ) ,.ICEIFA17 ( ICEIFA17 )
 ,.ICEIFA24 ( ICEIFA24 ) ,.ICEIFA16 ( ICEIFA16 ) ,.ICEIFA21 ( ICEIFA21 ) ,.ICEIFA13 ( ICEIFA13 ) ,.ICEIFA20 ( ICEIFA20 ) ,.ICEIFA12 ( ICEIFA12 )
 ,.ICEIFA11 ( ICEIFA11 ) ,.ICEIFA10 ( ICEIFA10 ) ,.ICEIFA9 ( ICEIFA9 ) ,.ICEIFA8 ( ICEIFA8 ) ,.ICEIFA7 ( ICEIFA7 ) ,.ICEIFA6 ( ICEIFA6 )
 ,.ICEIFA5 ( ICEIFA5 ) ,.ICEIFA4 ( ICEIFA4 ) ,.ICEIFA3 ( ICEIFA3 ) ,.ICEIFA2 ( ICEIFA2 ) ,.ICEIFA1 ( ICEIFA1 ) ,.ICEIFA0 ( ICEIFA0 )
 ,.ICEDI31 ( ICEDI31 ) ,.ICEDI23 ( ICEDI23 ) ,.ICEDI15 ( ICEDI15 ) ,.ICEDI30 ( ICEDI30 ) ,.ICEDI22 ( ICEDI22 ) ,.ICEDI14 ( ICEDI14 )
 ,.ICEDI29 ( ICEDI29 ) ,.ICEDI28 ( ICEDI28 ) ,.ICEDI27 ( ICEDI27 ) ,.ICEDI19 ( ICEDI19 ) ,.ICEDI26 ( ICEDI26 ) ,.ICEDI18 ( ICEDI18 )
 ,.ICEDI25 ( ICEDI25 ) ,.ICEDI17 ( ICEDI17 ) ,.ICEDI24 ( ICEDI24 ) ,.ICEDI16 ( ICEDI16 ) ,.ICEDI21 ( ICEDI21 ) ,.ICEDI13 ( ICEDI13 )
 ,.ICEDI20 ( ICEDI20 ) ,.ICEDI12 ( ICEDI12 ) ,.ICEDI11 ( ICEDI11 ) ,.ICEDI10 ( ICEDI10 ) ,.ICEDI9 ( ICEDI9 ) ,.ICEDI8 ( ICEDI8 )
 ,.ICEDI7 ( ICEDI7 ) ,.ICEDI6 ( ICEDI6 ) ,.ICEDI5 ( ICEDI5 ) ,.ICEDI4 ( ICEDI4 ) ,.ICEDI3 ( ICEDI3 ) ,.ICEDI2 ( ICEDI2 )
 ,.ICEDI1 ( ICEDI1 ) ,.ICEDI0 ( ICEDI0 ) ,.ICEWR ( ICEWR ) ,.EROMWAIT ( EROMWAIT ) ,.SVMOD ( SVMOD ) ,.SVMODF ( SVMODF )
 ,.ALT1 ( ALT1 ) ,.DW21 ( DW21 ) ,.DW13 ( DW13 ) ,.PREFIX ( PREFIX ) ,.SLFLASH ( SLFLASH ) ,.WAITFL2 ( WAITFL2 )
 ,.FLREAD ( FLREAD ) ,.PA19 ( PA19 ) ,.FCLK ( FCLK ) ,.PA18 ( PA18 ) ,.PA17 ( PA17 ) ,.PA16 ( PA16 )
 ,.PA15 ( PA15 ) ,.PA14 ( PA14 ) ,.PA13 ( PA13 ) ,.DW37 ( DW37 ) ,.DW29 ( DW29 ) ,.PA12 ( PA12 )
 ,.DW36 ( DW36 ) ,.DW28 ( DW28 ) ,.PA11 ( PA11 ) ,.DW35 ( DW35 ) ,.DW27 ( DW27 ) ,.DW19 ( DW19 )
 ,.PA10 ( PA10 ) ,.DW34 ( DW34 ) ,.DW26 ( DW26 ) ,.DW18 ( DW18 ) ,.PA9 ( PA9 ) ,.PA8 ( PA8 )
 ,.PA7 ( PA7 ) ,.PA6 ( PA6 ) ,.PA5 ( PA5 ) ,.DW9 ( DW9 ) ,.PA4 ( PA4 ) ,.DW8 ( DW8 )
 ,.PA3 ( PA3 ) ,.DIS ( DIS ) ,.DW7 ( DW7 ) ,.PA2 ( PA2 ) ,.DW6 ( DW6 ) ,.SLMEM ( SLMEM )
 ,.EXMA3 ( EXMA3 ) ,.RO137 ( RO137 ) ,.RO129 ( RO129 ) ,.EXMA2 ( EXMA2 ) ,.RO136 ( RO136 ) ,.RO128 ( RO128 )
 ,.EXMA1 ( EXMA1 ) ,.RO135 ( RO135 ) ,.RO127 ( RO127 ) ,.RO119 ( RO119 ) ,.EXMA0 ( EXMA0 ) ,.RO134 ( RO134 )
 ,.RO126 ( RO126 ) ,.RO118 ( RO118 ) ,.MA15 ( MA15 ) ,.MA14 ( MA14 ) ,.MA13 ( MA13 ) ,.MA12 ( MA12 )
 ,.BEU2 ( BEU2 ) ,.MA11 ( MA11 ) ,.BEU1 ( BEU1 ) ,.MA10 ( MA10 ) ,.BEU0 ( BEU0 ) ,.MA9 ( MA9 )
 ,.DW1 ( DW1 ) ,.MA8 ( MA8 ) ,.DW0 ( DW0 ) ,.MA7 ( MA7 ) ,.MA6 ( MA6 ) ,.MA5 ( MA5 )
 ,.MA4 ( MA4 ) ,.MA3 ( MA3 ) ,.MA2 ( MA2 ) ,.CER ( CER ) ,.MA1 ( MA1 ) ,.MA0 ( MA0 )
 ,.MDW15 ( MDW15 ) ,.MDW14 ( MDW14 ) ,.MDW13 ( MDW13 ) ,.MDW12 ( MDW12 ) ,.MDW11 ( MDW11 ) ,.MDW10 ( MDW10 )
 ,.MDW9 ( MDW9 ) ,.RO11 ( RO11 ) ,.RO03 ( RO03 ) ,.MDW8 ( MDW8 ) ,.RO10 ( RO10 ) ,.RO02 ( RO02 )
 ,.MDW7 ( MDW7 ) ,.RO01 ( RO01 ) ,.MDW6 ( MDW6 ) ,.RO00 ( RO00 ) ,.MDW5 ( MDW5 ) ,.MDW4 ( MDW4 )
 ,.MDW3 ( MDW3 ) ,.MDW2 ( MDW2 ) ,.MDW1 ( MDW1 ) ,.MDW0 ( MDW0 ) ,.EXCH ( EXCH ) ,.MEMMDR15 ( MEMMDR15 )
 ,.MEMMDR14 ( MEMMDR14 ) ,.MEMMDR13 ( MEMMDR13 ) ,.MEMMDR12 ( MEMMDR12 ) ,.MEMMDR11 ( MEMMDR11 ) ,.MEMMDR10 ( MEMMDR10 ) ,.MEMMDR9 ( MEMMDR9 )
 ,.MEMMDR8 ( MEMMDR8 ) ,.MEMMDR7 ( MEMMDR7 ) ,.MEMMDR6 ( MEMMDR6 ) ,.MEMMDR5 ( MEMMDR5 ) ,.MEMMDR4 ( MEMMDR4 ) ,.MEMMDR3 ( MEMMDR3 )
 ,.MEMMDR2 ( MEMMDR2 ) ,.MEMMDR1 ( MEMMDR1 ) ,.MEMMDR0 ( MEMMDR0 ) ,.CPUWR ( CPUWR ) ,.CPURD ( CPURD ) ,.RO020 ( RO020 )
 ,.RO012 ( RO012 ) ,.WDOP ( WDOP ) ,.FLMA15 ( FLMA15 ) ,.FLMA14 ( FLMA14 ) ,.FLMA13 ( FLMA13 ) ,.FLMA12 ( FLMA12 )
 ,.FLMA11 ( FLMA11 ) ,.FLMA10 ( FLMA10 ) ,.FLMA9 ( FLMA9 ) ,.FLMA8 ( FLMA8 ) ,.FLMA7 ( FLMA7 ) ,.FLMA6 ( FLMA6 )
 ,.FLMD0 ( FLMD0 ) ,.FLMA5 ( FLMA5 ) ,.FLMA4 ( FLMA4 ) ,.FLMA3 ( FLMA3 ) ,.FLMA2 ( FLMA2 ) ,.FLMA1 ( FLMA1 )
 ,.FLMA0 ( FLMA0 ) ,.SLBMEM ( SLBMEM ) ,.BRSAM ( BRSAM ) ,.FLSPMD ( FLSPMD ) ,.BTFLG ( BTFLG ) ,.TMSPMD ( TMSPMD )
 ,.TMBTSEL ( TMBTSEL ) ,.SWAP ( SWAP ) ,.ICETMSPMD ( ICETMSPMD ) ,.ICETMBTSEL ( ICETMBTSEL ) ,.RESB ( RESB ) ,.CLKSEL1 ( CLKSEL1 )
 ,.RDCLKP1 ( RDCLKP1 ) ,.CE0 ( CE0 ) ,.CE1 ( CE1 ) ,.EXA ( EXA ) ,.A19 ( A19 ) ,.A18 ( A18 )
 ,.A17 ( A17 ) ,.A16 ( A16 ) ,.A15 ( A15 ) ,.A14 ( A14 ) ,.A13 ( A13 ) ,.A12 ( A12 )
 ,.A11 ( A11 ) ,.A10 ( A10 ) ,.A9 ( A9 ) ,.A8 ( A8 ) ,.A7 ( A7 ) ,.A6 ( A6 )
 ,.A5 ( A5 ) ,.A4 ( A4 ) ,.A3 ( A3 ) ,.A2 ( A2 ) ,.RO133 ( RO133 ) ,.RO125 ( RO125 )
 ,.RO117 ( RO117 ) ,.RO037 ( RO037 ) ,.RO029 ( RO029 ) ,.RO132 ( RO132 ) ,.RO124 ( RO124 ) ,.RO116 ( RO116 )
 ,.RO036 ( RO036 ) ,.RO028 ( RO028 ) ,.RO131 ( RO131 ) ,.RO123 ( RO123 ) ,.RO115 ( RO115 ) ,.RO035 ( RO035 )
 ,.RO027 ( RO027 ) ,.RO019 ( RO019 ) ,.RO130 ( RO130 ) ,.RO122 ( RO122 ) ,.RO114 ( RO114 ) ,.RO034 ( RO034 )
 ,.RO026 ( RO026 ) ,.RO018 ( RO018 ) ,.RO121 ( RO121 ) ,.RO113 ( RO113 ) ,.RO033 ( RO033 ) ,.RO025 ( RO025 )
 ,.RO017 ( RO017 ) ,.RO120 ( RO120 ) ,.RO112 ( RO112 ) ,.RO032 ( RO032 ) ,.RO024 ( RO024 ) ,.RO016 ( RO016 )
 ,.RO111 ( RO111 ) ,.RO031 ( RO031 ) ,.RO023 ( RO023 ) ,.RO015 ( RO015 ) ,.RO110 ( RO110 ) ,.RO030 ( RO030 )
 ,.RO022 ( RO022 ) ,.RO014 ( RO014 ) ,.RO19 ( RO19 ) ,.RO18 ( RO18 ) ,.RO17 ( RO17 ) ,.RO09 ( RO09 )
 ,.RO16 ( RO16 ) ,.RO08 ( RO08 ) ,.RO15 ( RO15 ) ,.RO07 ( RO07 ) ,.RO14 ( RO14 ) ,.RO06 ( RO06 )
 ,.RO13 ( RO13 ) ,.RO05 ( RO05 ) ,.RO12 ( RO12 ) ,.RO04 ( RO04 ) ,.RO021 ( RO021 ) ,.RO013 ( RO013 )
 ,.RO011 ( RO011 ) ,.RO010 ( RO010 ) ,.SELRO1 ( SELRO1 ) ,.CIBPID31 ( CIBPID31 ) ,.CIBPID23 ( CIBPID23 ) ,.CIBPID15 ( CIBPID15 )
 ,.CIBPID30 ( CIBPID30 ) ,.CIBPID22 ( CIBPID22 ) ,.CIBPID14 ( CIBPID14 ) ,.CIBPID29 ( CIBPID29 ) ,.CIBPID28 ( CIBPID28 ) ,.CIBPID27 ( CIBPID27 )
 ,.CIBPID19 ( CIBPID19 ) ,.CIBPID26 ( CIBPID26 ) ,.CIBPID18 ( CIBPID18 ) ,.CIBPID25 ( CIBPID25 ) ,.CIBPID17 ( CIBPID17 ) ,.CIBPID24 ( CIBPID24 )
 ,.CIBPID16 ( CIBPID16 ) ,.CIBPID21 ( CIBPID21 ) ,.CIBPID13 ( CIBPID13 ) ,.CIBPID20 ( CIBPID20 ) ,.CIBPID12 ( CIBPID12 ) ,.CIBPID11 ( CIBPID11 )
 ,.CIBPID10 ( CIBPID10 ) ,.CIBPID9 ( CIBPID9 ) ,.CIBPID8 ( CIBPID8 ) ,.CIBPID7 ( CIBPID7 ) ,.CIBPID6 ( CIBPID6 ) ,.CIBPID5 ( CIBPID5 )
 ,.CIBPID4 ( CIBPID4 ) ,.CIBPID3 ( CIBPID3 ) ,.CIBPID2 ( CIBPID2 ) ,.CIBPID1 ( CIBPID1 ) ,.CIBPID0 ( CIBPID0 ) ,.CPUPID31 ( CPUPID31 )
 ,.CPUPID23 ( CPUPID23 ) ,.CPUPID15 ( CPUPID15 ) ,.CPUPID30 ( CPUPID30 ) ,.CPUPID22 ( CPUPID22 ) ,.CPUPID14 ( CPUPID14 ) ,.CPUPID29 ( CPUPID29 )
 ,.CPUPID28 ( CPUPID28 ) ,.CPUPID27 ( CPUPID27 ) ,.CPUPID19 ( CPUPID19 ) ,.CPUPID26 ( CPUPID26 ) ,.CPUPID18 ( CPUPID18 ) ,.CPUPID25 ( CPUPID25 )
 ,.CPUPID17 ( CPUPID17 ) ,.CPUPID24 ( CPUPID24 ) ,.CPUPID16 ( CPUPID16 ) ,.CPUPID21 ( CPUPID21 ) ,.CPUPID13 ( CPUPID13 ) ,.CPUPID20 ( CPUPID20 )
 ,.CPUPID12 ( CPUPID12 ) ,.CPUPID11 ( CPUPID11 ) ,.CPUPID10 ( CPUPID10 ) ,.CPUPID9 ( CPUPID9 ) ,.CPUPID8 ( CPUPID8 ) ,.CPUPID7 ( CPUPID7 )
 ,.CPUPID6 ( CPUPID6 ) ,.CPUPID5 ( CPUPID5 ) ,.CPUPID4 ( CPUPID4 ) ,.CPUPID3 ( CPUPID3 ) ,.CPUPID2 ( CPUPID2 ) ,.CPUPID1 ( CPUPID1 )
 ,.CPUPID0 ( CPUPID0 ) ,.WWR ( WWR ) ,.SER ( SER ) ,.MRG00 ( MRG00 ) ,.MRG01 ( MRG01 ) ,.MRG10 ( MRG10 )
 ,.MRG11 ( MRG11 ) ,.MRG12 ( MRG12 ) ,.READ ( READ ) ,.PROGI ( PROGI ) ,.WED ( WED ) ,.BFA ( BFA )
 ,.DW33 ( DW33 ) ,.DW25 ( DW25 ) ,.DW17 ( DW17 ) ,.DW32 ( DW32 ) ,.DW24 ( DW24 ) ,.DW16 ( DW16 )
 ,.DW31 ( DW31 ) ,.DW23 ( DW23 ) ,.DW15 ( DW15 ) ,.DW30 ( DW30 ) ,.DW22 ( DW22 ) ,.DW14 ( DW14 )
 ,.DW20 ( DW20 ) ,.DW12 ( DW12 ) ,.DW11 ( DW11 ) ,.DW10 ( DW10 ) ,.DW5 ( DW5 ) ,.DW4 ( DW4 )
 ,.DW3 ( DW3 ) ,.DW2 ( DW2 ) ,.ICENOECC ( ICENOECC ) ,.MAAOUT ( MAAOUT ) ,.SELFMODE ( SELFMODE ) ,.SELFMODEDBG ( SELFMODEDBG )
 ,.FAILMK12 ( FAILMK12 ) ,.BRKFAIL12 ( BRKFAIL12 ) ,.BFBRKPID31 ( BFBRKPID31 ) ,.BFBRKPID23 ( BFBRKPID23 ) ,.BFBRKPID15 ( BFBRKPID15 ) ,.BFBRKPID30 ( BFBRKPID30 )
 ,.BFBRKPID22 ( BFBRKPID22 ) ,.BFBRKPID14 ( BFBRKPID14 ) ,.BFBRKPID29 ( BFBRKPID29 ) ,.BFBRKPID28 ( BFBRKPID28 ) ,.BFBRKPID27 ( BFBRKPID27 ) ,.BFBRKPID19 ( BFBRKPID19 )
 ,.BFBRKPID26 ( BFBRKPID26 ) ,.BFBRKPID18 ( BFBRKPID18 ) ,.BFBRKPID25 ( BFBRKPID25 ) ,.BFBRKPID17 ( BFBRKPID17 ) ,.BFBRKPID24 ( BFBRKPID24 ) ,.BFBRKPID16 ( BFBRKPID16 )
 ,.BFBRKPID21 ( BFBRKPID21 ) ,.BFBRKPID13 ( BFBRKPID13 ) ,.BFBRKPID20 ( BFBRKPID20 ) ,.BFBRKPID12 ( BFBRKPID12 ) ,.BFBRKPID11 ( BFBRKPID11 ) ,.BFBRKPID10 ( BFBRKPID10 )
 ,.BFBRKPID9 ( BFBRKPID9 ) ,.BFBRKPID8 ( BFBRKPID8 ) ,.BFBRKPID7 ( BFBRKPID7 ) ,.BFBRKPID6 ( BFBRKPID6 ) ,.BFBRKPID5 ( BFBRKPID5 ) ,.BFBRKPID4 ( BFBRKPID4 )
 ,.BFBRKPID3 ( BFBRKPID3 ) ,.BFBRKPID2 ( BFBRKPID2 ) ,.BFBRKPID1 ( BFBRKPID1 ) ,.BFBRKPID0 ( BFBRKPID0 ) ,.GDRAMWR ( GDRAMWR ) ,.SYSRSOUTB ( SYSRSOUTB )
 ,.BASECK ( BASECK ) ,.EMEMRAMCLK ( EMEMRAMCLK )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/bforebreak.v
  BFOREBREAK bforebreak (
   .ICEDO31 ( ICEDOD31 ) ,.ICEDO23 ( ICEDOD23 ) ,.ICEDO15 ( ICEDOD15 ) ,.ICEDO30 ( ICEDOD30 ) ,.ICEDO22 ( ICEDOD22 ) ,.ICEDO14 ( ICEDOD14 ) ,.ICEDO29 ( ICEDOD29 )
 ,.ICEDO28 ( ICEDOD28 ) ,.ICEDO27 ( ICEDOD27 ) ,.ICEDO19 ( ICEDOD19 ) ,.ICEDO26 ( ICEDOD26 ) ,.ICEDO18 ( ICEDOD18 ) ,.ICEDO25 ( ICEDOD25 )
 ,.ICEDO17 ( ICEDOD17 ) ,.ICEDO24 ( ICEDOD24 ) ,.ICEDO16 ( ICEDOD16 ) ,.ICEDO21 ( ICEDOD21 ) ,.ICEDO13 ( ICEDOD13 ) ,.ICEDO20 ( ICEDOD20 )
 ,.ICEDO12 ( ICEDOD12 ) ,.ICEDO11 ( ICEDOD11 ) ,.ICEDO10 ( ICEDOD10 ) ,.ICEDO9 ( ICEDOD9 ) ,.ICEDO8 ( ICEDOD8 ) ,.ICEDO7 ( ICEDOD7 )
 ,.ICEDO6 ( ICEDOD6 ) ,.ICEDO5 ( ICEDOD5 ) ,.ICEDO4 ( ICEDOD4 ) ,.ICEDO3 ( ICEDOD3 ) ,.ICEDO2 ( ICEDOD2 ) ,.ICEDO1 ( ICEDOD1 )
 ,.ICEDO0 ( ICEDOD0 ) ,.ICEIFA31 ( ICEIFA31 ) ,.ICEIFA23 ( ICEIFA23 ) ,.ICEIFA15 ( ICEIFA15 ) ,.ICEIFA30 ( ICEIFA30 ) ,.ICEIFA22 ( ICEIFA22 )
 ,.ICEIFA14 ( ICEIFA14 ) ,.ICEIFA29 ( ICEIFA29 ) ,.ICEIFA28 ( ICEIFA28 ) ,.ICEIFA27 ( ICEIFA27 ) ,.ICEIFA19 ( ICEIFA19 ) ,.ICEIFA26 ( ICEIFA26 )
 ,.ICEIFA18 ( ICEIFA18 ) ,.ICEIFA25 ( ICEIFA25 ) ,.ICEIFA17 ( ICEIFA17 ) ,.ICEIFA24 ( ICEIFA24 ) ,.ICEIFA16 ( ICEIFA16 ) ,.ICEIFA21 ( ICEIFA21 )
 ,.ICEIFA13 ( ICEIFA13 ) ,.ICEIFA20 ( ICEIFA20 ) ,.ICEIFA12 ( ICEIFA12 ) ,.ICEIFA11 ( ICEIFA11 ) ,.ICEIFA10 ( ICEIFA10 ) ,.ICEIFA9 ( ICEIFA9 )
 ,.ICEIFA8 ( ICEIFA8 ) ,.ICEIFA7 ( ICEIFA7 ) ,.ICEIFA6 ( ICEIFA6 ) ,.ICEIFA5 ( ICEIFA5 ) ,.ICEIFA4 ( ICEIFA4 ) ,.ICEIFA3 ( ICEIFA3 )
 ,.ICEIFA2 ( ICEIFA2 ) ,.ICEIFA1 ( ICEIFA1 ) ,.ICEIFA0 ( ICEIFA0 ) ,.ICEDI31 ( ICEDI31 ) ,.ICEDI23 ( ICEDI23 ) ,.ICEDI15 ( ICEDI15 )
 ,.ICEDI30 ( ICEDI30 ) ,.ICEDI22 ( ICEDI22 ) ,.ICEDI14 ( ICEDI14 ) ,.ICEDI29 ( ICEDI29 ) ,.ICEDI28 ( ICEDI28 ) ,.ICEDI27 ( ICEDI27 )
 ,.ICEDI19 ( ICEDI19 ) ,.ICEDI26 ( ICEDI26 ) ,.ICEDI18 ( ICEDI18 ) ,.ICEDI25 ( ICEDI25 ) ,.ICEDI17 ( ICEDI17 ) ,.ICEDI24 ( ICEDI24 )
 ,.ICEDI16 ( ICEDI16 ) ,.ICEDI21 ( ICEDI21 ) ,.ICEDI13 ( ICEDI13 ) ,.ICEDI20 ( ICEDI20 ) ,.ICEDI12 ( ICEDI12 ) ,.ICEDI11 ( ICEDI11 )
 ,.ICEDI10 ( ICEDI10 ) ,.ICEDI9 ( ICEDI9 ) ,.ICEDI8 ( ICEDI8 ) ,.ICEDI7 ( ICEDI7 ) ,.ICEDI6 ( ICEDI6 ) ,.ICEDI5 ( ICEDI5 )
 ,.ICEDI4 ( ICEDI4 ) ,.ICEDI3 ( ICEDI3 ) ,.ICEDI2 ( ICEDI2 ) ,.ICEDI1 ( ICEDI1 ) ,.ICEDI0 ( ICEDI0 ) ,.ICEWR ( ICEWR )
 ,.PA19 ( PA19 ) ,.PA18 ( PA18 ) ,.PA17 ( PA17 ) ,.PA16 ( PA16 ) ,.PA15 ( PA15 ) ,.PA14 ( PA14 )
 ,.PA13 ( PA13 ) ,.PA12 ( PA12 ) ,.PA11 ( PA11 ) ,.PA10 ( PA10 ) ,.PA9 ( PA9 ) ,.PA8 ( PA8 )
 ,.PA7 ( PA7 ) ,.PA6 ( PA6 ) ,.PA5 ( PA5 ) ,.PA4 ( PA4 ) ,.PA3 ( PA3 ) ,.PA2 ( PA2 )
 ,.BFBRKPID31 ( BFBRKPID31 ) ,.BFBRKPID23 ( BFBRKPID23 ) ,.BFBRKPID15 ( BFBRKPID15 ) ,.BFBRKPID30 ( BFBRKPID30 ) ,.BFBRKPID22 ( BFBRKPID22 ) ,.BFBRKPID14 ( BFBRKPID14 )
 ,.BFBRKPID29 ( BFBRKPID29 ) ,.BFBRKPID28 ( BFBRKPID28 ) ,.BFBRKPID27 ( BFBRKPID27 ) ,.BFBRKPID19 ( BFBRKPID19 ) ,.BFBRKPID26 ( BFBRKPID26 ) ,.BFBRKPID18 ( BFBRKPID18 )
 ,.BFBRKPID25 ( BFBRKPID25 ) ,.BFBRKPID17 ( BFBRKPID17 ) ,.BFBRKPID24 ( BFBRKPID24 ) ,.BFBRKPID16 ( BFBRKPID16 ) ,.BFBRKPID21 ( BFBRKPID21 ) ,.BFBRKPID13 ( BFBRKPID13 )
 ,.BFBRKPID20 ( BFBRKPID20 ) ,.BFBRKPID12 ( BFBRKPID12 ) ,.BFBRKPID11 ( BFBRKPID11 ) ,.BFBRKPID10 ( BFBRKPID10 ) ,.BFBRKPID9 ( BFBRKPID9 ) ,.BFBRKPID8 ( BFBRKPID8 )
 ,.BFBRKPID7 ( BFBRKPID7 ) ,.BFBRKPID6 ( BFBRKPID6 ) ,.BFBRKPID5 ( BFBRKPID5 ) ,.BFBRKPID4 ( BFBRKPID4 ) ,.BFBRKPID3 ( BFBRKPID3 ) ,.BFBRKPID2 ( BFBRKPID2 )
 ,.BFBRKPID1 ( BFBRKPID1 ) ,.BFBRKPID0 ( BFBRKPID0 ) ,.BFBRKSEL ( BFBRKSEL ) ,.SYSRSOUTB ( SYSRSOUTB ) ,.BASECK ( BASECK ) ,.FLREAD ( FLREAD )
 ,.SVMODF ( SVMODF ) ,.PCWAITF ( PCWAITF )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/host_interface.v
  HOST_INTERFACE host_interface (
   .ICESYSRES_B ( EICESYSRES_B ) ,.CLK60MHZ ( CLK30MHZ_GB ) ,.EROMWAIT ( WAITOR ) ,.CPURESETB ( CPURSOUTB ) ,.ES3 ( EXMA3 ) ,.MA7 ( MA7 ) ,.ES2 ( EXMA2 )
 ,.MA6 ( MA6 ) ,.ES1 ( EXMA1 ) ,.MA5 ( MA5 ) ,.ES0 ( EXMA0 ) ,.MA4 ( MA4 ) ,.MDR15 ( HOSTIFMDR15 )
 ,.MDR14 ( HOSTIFMDR14 ) ,.MDR13 ( HOSTIFMDR13 ) ,.MDR12 ( HOSTIFMDR12 ) ,.MDR11 ( HOSTIFMDR11 ) ,.MDR10 ( HOSTIFMDR10 ) ,.MDR9 ( HOSTIFMDR9 )
 ,.MDR8 ( HOSTIFMDR8 ) ,.MDR7 ( HOSTIFMDR7 ) ,.MDR6 ( HOSTIFMDR6 ) ,.MDR5 ( HOSTIFMDR5 ) ,.MDR4 ( HOSTIFMDR4 ) ,.MDR3 ( HOSTIFMDR3 )
 ,.MDR2 ( HOSTIFMDR2 ) ,.MDR1 ( HOSTIFMDR1 ) ,.MDR0 ( HOSTIFMDR0 ) ,.USBCLK ( USBCLK ) ,.USBA21 ( USBA21 ) ,.USBA20 ( USBA20 )
 ,.USBA19 ( USBA19 ) ,.USBA4 ( USBA4 ) ,.USBA3 ( USBA3 ) ,.USBA2 ( USBA2 ) ,.USBA1 ( USBA1 ) ,.USBD15 ( USBD15 )
 ,.USBD14 ( USBD14 ) ,.USBD13 ( USBD13 ) ,.USBD12 ( USBD12 ) ,.USBD11 ( USBD11 ) ,.USBD10 ( USBD10 ) ,.USBD9 ( USBD9 )
 ,.USBD8 ( USBD8 ) ,.USBD7 ( USBD7 ) ,.USBD6 ( USBD6 ) ,.USBD5 ( USBD5 ) ,.USBD4 ( USBD4 ) ,.USBD3 ( USBD3 )
 ,.USBD2 ( USBD2 ) ,.USBD1 ( USBD1 ) ,.USBD0 ( USBD0 ) ,.USBRD_B ( USBRD_B ) ,.USBWR0_B ( USBWR0_B ) ,.USBWAIT_B ( USBWAIT_B )
 ,.ICEIFA31 ( ICEIFA31 ) ,.ICEIFA23 ( ICEIFA23 ) ,.ICEIFA15 ( ICEIFA15 ) ,.ICEDOB27 ( ICEDOB27 ) ,.ICEDOB19 ( ICEDOB19 ) ,.ICEDOC31 ( ICEDOC31 )
 ,.ICEDOC23 ( ICEDOC23 ) ,.ICEDOC15 ( ICEDOC15 ) ,.ICEDOD11 ( ICEDOD11 ) ,.ICEIFA30 ( ICEIFA30 ) ,.ICEIFA22 ( ICEIFA22 ) ,.ICEIFA14 ( ICEIFA14 )
 ,.ICEDOB26 ( ICEDOB26 ) ,.ICEDOB18 ( ICEDOB18 ) ,.ICEDOC30 ( ICEDOC30 ) ,.ICEDOC22 ( ICEDOC22 ) ,.ICEDOC14 ( ICEDOC14 ) ,.ICEDOD10 ( ICEDOD10 )
 ,.ICEIFA29 ( ICEIFA29 ) ,.ICEDOC29 ( ICEDOC29 ) ,.ICEDOD25 ( ICEDOD25 ) ,.ICEDOD17 ( ICEDOD17 ) ,.ICEDOE21 ( ICEDOE21 ) ,.ICEDOE13 ( ICEDOE13 )
 ,.ICEIFA28 ( ICEIFA28 ) ,.ICEDOC28 ( ICEDOC28 ) ,.ICEDOD24 ( ICEDOD24 ) ,.ICEDOD16 ( ICEDOD16 ) ,.ICEDOE20 ( ICEDOE20 ) ,.ICEDOE12 ( ICEDOE12 )
 ,.ICEIFA27 ( ICEIFA27 ) ,.ICEIFA19 ( ICEIFA19 ) ,.ICEDOC27 ( ICEDOC27 ) ,.ICEDOC19 ( ICEDOC19 ) ,.ICEDOD31 ( ICEDOD31 ) ,.ICEDOD23 ( ICEDOD23 )
 ,.ICEDOD15 ( ICEDOD15 ) ,.ICEDOE11 ( ICEDOE11 ) ,.ICEIFA26 ( ICEIFA26 ) ,.ICEIFA18 ( ICEIFA18 ) ,.ICEDOC26 ( ICEDOC26 ) ,.ICEDOC18 ( ICEDOC18 )
 ,.ICEDOD30 ( ICEDOD30 ) ,.ICEDOD22 ( ICEDOD22 ) ,.ICEDOD14 ( ICEDOD14 ) ,.ICEDOE10 ( ICEDOE10 ) ,.ICEIFA25 ( ICEIFA25 ) ,.ICEIFA17 ( ICEIFA17 )
 ,.ICEDOB29 ( ICEDOB29 ) ,.ICEDOC25 ( ICEDOC25 ) ,.ICEDOC17 ( ICEDOC17 ) ,.ICEDOD21 ( ICEDOD21 ) ,.ICEDOD13 ( ICEDOD13 ) ,.ICEIFA24 ( ICEIFA24 )
 ,.ICEIFA16 ( ICEIFA16 ) ,.ICEDOB28 ( ICEDOB28 ) ,.ICEDOC24 ( ICEDOC24 ) ,.ICEDOC16 ( ICEDOC16 ) ,.ICEDOD20 ( ICEDOD20 ) ,.ICEDOD12 ( ICEDOD12 )
 ,.ICEIFA21 ( ICEIFA21 ) ,.ICEIFA13 ( ICEIFA13 ) ,.ICEDOA29 ( ICEDOA29 ) ,.ICEDOB25 ( ICEDOB25 ) ,.ICEDOB17 ( ICEDOB17 ) ,.ICEDOC21 ( ICEDOC21 )
 ,.ICEDOC13 ( ICEDOC13 ) ,.ICEIFA20 ( ICEIFA20 ) ,.ICEIFA12 ( ICEIFA12 ) ,.ICEDOA28 ( ICEDOA28 ) ,.ICEDOB24 ( ICEDOB24 ) ,.ICEDOB16 ( ICEDOB16 )
 ,.ICEDOC20 ( ICEDOC20 ) ,.ICEDOC12 ( ICEDOC12 ) ,.ICEIFA11 ( ICEIFA11 ) ,.ICEDOA27 ( ICEDOA27 ) ,.ICEDOA19 ( ICEDOA19 ) ,.ICEDOB31 ( ICEDOB31 )
 ,.ICEDOB23 ( ICEDOB23 ) ,.ICEDOB15 ( ICEDOB15 ) ,.ICEDOC11 ( ICEDOC11 ) ,.ICEIFA10 ( ICEIFA10 ) ,.ICEDOA26 ( ICEDOA26 ) ,.ICEDOA18 ( ICEDOA18 )
 ,.ICEDOB30 ( ICEDOB30 ) ,.ICEDOB22 ( ICEDOB22 ) ,.ICEDOB14 ( ICEDOB14 ) ,.ICEDOC10 ( ICEDOC10 ) ,.ICEIFA9 ( ICEIFA9 ) ,.ICEDOC9 ( ICEDOC9 )
 ,.ICEDOD7 ( ICEDOD7 ) ,.ICEDOE5 ( ICEDOE5 ) ,.ICEDOF3 ( ICEDOF3 ) ,.ICEDOG1 ( ICEDOG1 ) ,.ICEIFA8 ( ICEIFA8 ) ,.ICEDOC8 ( ICEDOC8 )
 ,.ICEDOD6 ( ICEDOD6 ) ,.ICEDOE4 ( ICEDOE4 ) ,.ICEDOF2 ( ICEDOF2 ) ,.ICEDOG0 ( ICEDOG0 ) ,.ICEIFA7 ( ICEIFA7 ) ,.ICEDOB9 ( ICEDOB9 )
 ,.ICEDOC7 ( ICEDOC7 ) ,.ICEDOD5 ( ICEDOD5 ) ,.ICEDOE3 ( ICEDOE3 ) ,.ICEDOF1 ( ICEDOF1 ) ,.ICEIFA6 ( ICEIFA6 ) ,.ICEDOB8 ( ICEDOB8 )
 ,.ICEDOC6 ( ICEDOC6 ) ,.ICEDOD4 ( ICEDOD4 ) ,.ICEDOE2 ( ICEDOE2 ) ,.ICEDOF0 ( ICEDOF0 ) ,.ICEIFA5 ( ICEIFA5 ) ,.ICEDOA9 ( ICEDOA9 )
 ,.ICEDOB7 ( ICEDOB7 ) ,.ICEDOC5 ( ICEDOC5 ) ,.ICEDOD3 ( ICEDOD3 ) ,.ICEDOE1 ( ICEDOE1 ) ,.ICEIFA4 ( ICEIFA4 ) ,.ICEDOA8 ( ICEDOA8 )
 ,.ICEDOB6 ( ICEDOB6 ) ,.ICEDOC4 ( ICEDOC4 ) ,.ICEDOD2 ( ICEDOD2 ) ,.ICEDOE0 ( ICEDOE0 ) ,.ICEIFA3 ( ICEIFA3 ) ,.ICEDOA7 ( ICEDOA7 )
 ,.ICEDOB5 ( ICEDOB5 ) ,.ICEDOC3 ( ICEDOC3 ) ,.ICEDOD1 ( ICEDOD1 ) ,.ICEIFA2 ( ICEIFA2 ) ,.ICEDOA6 ( ICEDOA6 ) ,.ICEDOB4 ( ICEDOB4 )
 ,.ICEDOC2 ( ICEDOC2 ) ,.ICEDOD0 ( ICEDOD0 ) ,.ICEIFA1 ( ICEIFA1 ) ,.ICEDOA5 ( ICEDOA5 ) ,.ICEDOB3 ( ICEDOB3 ) ,.ICEDOC1 ( ICEDOC1 )
 ,.ICEIFA0 ( ICEIFA0 ) ,.ICEDOA4 ( ICEDOA4 ) ,.ICEDOB2 ( ICEDOB2 ) ,.ICEDOC0 ( ICEDOC0 ) ,.ICEDOA31 ( ICEDOA31 ) ,.ICEDOA23 ( ICEDOA23 )
 ,.ICEDOA15 ( ICEDOA15 ) ,.ICEDOB11 ( ICEDOB11 ) ,.ICEDOA30 ( ICEDOA30 ) ,.ICEDOA22 ( ICEDOA22 ) ,.ICEDOA14 ( ICEDOA14 ) ,.ICEDOB10 ( ICEDOB10 )
 ,.ICEDOA25 ( ICEDOA25 ) ,.ICEDOA17 ( ICEDOA17 ) ,.ICEDOB21 ( ICEDOB21 ) ,.ICEDOB13 ( ICEDOB13 ) ,.ICEDOA24 ( ICEDOA24 ) ,.ICEDOA16 ( ICEDOA16 )
 ,.ICEDOB20 ( ICEDOB20 ) ,.ICEDOB12 ( ICEDOB12 ) ,.ICEDOA21 ( ICEDOA21 ) ,.ICEDOA13 ( ICEDOA13 ) ,.ICEDOA20 ( ICEDOA20 ) ,.ICEDOA12 ( ICEDOA12 )
 ,.ICEDOA11 ( ICEDOA11 ) ,.ICEDOA10 ( ICEDOA10 ) ,.ICEDOA3 ( ICEDOA3 ) ,.ICEDOB1 ( ICEDOB1 ) ,.ICEDOA2 ( ICEDOA2 ) ,.ICEDOB0 ( ICEDOB0 )
 ,.ICEDOA1 ( ICEDOA1 ) ,.ICEDOA0 ( ICEDOA0 ) ,.ICEDOD29 ( ICEDOD29 ) ,.ICEDOE25 ( ICEDOE25 ) ,.ICEDOE17 ( ICEDOE17 ) ,.ICEDOF21 ( ICEDOF21 )
 ,.ICEDOF13 ( ICEDOF13 ) ,.ICEDOD28 ( ICEDOD28 ) ,.ICEDOE24 ( ICEDOE24 ) ,.ICEDOE16 ( ICEDOE16 ) ,.ICEDOF20 ( ICEDOF20 ) ,.ICEDOF12 ( ICEDOF12 )
 ,.ICEDOD27 ( ICEDOD27 ) ,.ICEDOD19 ( ICEDOD19 ) ,.ICEDOE31 ( ICEDOE31 ) ,.ICEDOE23 ( ICEDOE23 ) ,.ICEDOE15 ( ICEDOE15 ) ,.ICEDOF11 ( ICEDOF11 )
 ,.ICEDOD26 ( ICEDOD26 ) ,.ICEDOD18 ( ICEDOD18 ) ,.ICEDOE30 ( ICEDOE30 ) ,.ICEDOE22 ( ICEDOE22 ) ,.ICEDOE14 ( ICEDOE14 ) ,.ICEDOF10 ( ICEDOF10 )
 ,.ICEDOD9 ( ICEDOD9 ) ,.ICEDOE7 ( ICEDOE7 ) ,.ICEDOF5 ( ICEDOF5 ) ,.ICEDOG3 ( ICEDOG3 ) ,.ICEDOH1 ( ICEDOH1 ) ,.ICEDOD8 ( ICEDOD8 )
 ,.ICEDOE6 ( ICEDOE6 ) ,.ICEDOF4 ( ICEDOF4 ) ,.ICEDOG2 ( ICEDOG2 ) ,.ICEDOH0 ( ICEDOH0 ) ,.ICEDOE29 ( ICEDOE29 ) ,.ICEDOF25 ( ICEDOF25 )
 ,.ICEDOF17 ( ICEDOF17 ) ,.ICEDOG21 ( ICEDOG21 ) ,.ICEDOG13 ( ICEDOG13 ) ,.ICEDOE28 ( ICEDOE28 ) ,.ICEDOF24 ( ICEDOF24 ) ,.ICEDOF16 ( ICEDOF16 )
 ,.ICEDOG20 ( ICEDOG20 ) ,.ICEDOG12 ( ICEDOG12 ) ,.ICEDOE27 ( ICEDOE27 ) ,.ICEDOE19 ( ICEDOE19 ) ,.ICEDOF31 ( ICEDOF31 ) ,.ICEDOF23 ( ICEDOF23 )
 ,.ICEDOF15 ( ICEDOF15 ) ,.ICEDOG11 ( ICEDOG11 ) ,.ICEDOE26 ( ICEDOE26 ) ,.ICEDOE18 ( ICEDOE18 ) ,.ICEDOF30 ( ICEDOF30 ) ,.ICEDOF22 ( ICEDOF22 )
 ,.ICEDOF14 ( ICEDOF14 ) ,.ICEDOG10 ( ICEDOG10 ) ,.ICEDOE9 ( ICEDOE9 ) ,.ICEDOF7 ( ICEDOF7 ) ,.ICEDOG5 ( ICEDOG5 ) ,.ICEDOH3 ( ICEDOH3 )
 ,.ICEDOE8 ( ICEDOE8 ) ,.ICEDOF6 ( ICEDOF6 ) ,.ICEDOG4 ( ICEDOG4 ) ,.ICEDOH2 ( ICEDOH2 ) ,.ICEDOF29 ( ICEDOF29 ) ,.ICEDOG25 ( ICEDOG25 )
 ,.ICEDOG17 ( ICEDOG17 ) ,.ICEDOH21 ( ICEDOH21 ) ,.ICEDOH13 ( ICEDOH13 ) ,.ICEDOF28 ( ICEDOF28 ) ,.ICEDOG24 ( ICEDOG24 ) ,.ICEDOG16 ( ICEDOG16 )
 ,.ICEDOH20 ( ICEDOH20 ) ,.ICEDOH12 ( ICEDOH12 ) ,.ICEDOF27 ( ICEDOF27 ) ,.ICEDOF19 ( ICEDOF19 ) ,.ICEDOG31 ( ICEDOG31 ) ,.ICEDOG23 ( ICEDOG23 )
 ,.ICEDOG15 ( ICEDOG15 ) ,.ICEDOH11 ( ICEDOH11 ) ,.ICEDOF26 ( ICEDOF26 ) ,.ICEDOF18 ( ICEDOF18 ) ,.ICEDOG30 ( ICEDOG30 ) ,.ICEDOG22 ( ICEDOG22 )
 ,.ICEDOG14 ( ICEDOG14 ) ,.ICEDOH10 ( ICEDOH10 ) ,.ICEDOF9 ( ICEDOF9 ) ,.ICEDOG7 ( ICEDOG7 ) ,.ICEDOH5 ( ICEDOH5 ) ,.ICEDOJ1 ( ICEDOJ1 )
 ,.ICEDOF8 ( ICEDOF8 ) ,.ICEDOG6 ( ICEDOG6 ) ,.ICEDOH4 ( ICEDOH4 ) ,.ICEDOJ0 ( ICEDOJ0 ) ,.ICEDOG29 ( ICEDOG29 ) ,.ICEDOH25 ( ICEDOH25 )
 ,.ICEDOH17 ( ICEDOH17 ) ,.ICEDOG28 ( ICEDOG28 ) ,.ICEDOH24 ( ICEDOH24 ) ,.ICEDOH16 ( ICEDOH16 ) ,.ICEDOG27 ( ICEDOG27 ) ,.ICEDOG19 ( ICEDOG19 )
 ,.ICEDOH31 ( ICEDOH31 ) ,.ICEDOH23 ( ICEDOH23 ) ,.ICEDOH15 ( ICEDOH15 ) ,.ICEDOG26 ( ICEDOG26 ) ,.ICEDOG18 ( ICEDOG18 ) ,.ICEDOH30 ( ICEDOH30 )
 ,.ICEDOH22 ( ICEDOH22 ) ,.ICEDOH14 ( ICEDOH14 ) ,.ICEDOG9 ( ICEDOG9 ) ,.ICEDOH7 ( ICEDOH7 ) ,.ICEDOJ3 ( ICEDOJ3 ) ,.ICEDOK1 ( ICEDOK1 )
 ,.ICEDOG8 ( ICEDOG8 ) ,.ICEDOH6 ( ICEDOH6 ) ,.ICEDOJ2 ( ICEDOJ2 ) ,.ICEDOK0 ( ICEDOK0 ) ,.ICEDOH29 ( ICEDOH29 ) ,.ICEDOJ21 ( ICEDOJ21 )
 ,.ICEDOJ13 ( ICEDOJ13 ) ,.ICEDOH28 ( ICEDOH28 ) ,.ICEDOJ20 ( ICEDOJ20 ) ,.ICEDOJ12 ( ICEDOJ12 ) ,.ICEDOH27 ( ICEDOH27 ) ,.ICEDOH19 ( ICEDOH19 )
 ,.ICEDOJ11 ( ICEDOJ11 ) ,.ICEDOH26 ( ICEDOH26 ) ,.ICEDOH18 ( ICEDOH18 ) ,.ICEDOJ10 ( ICEDOJ10 ) ,.ICEDOH9 ( ICEDOH9 ) ,.ICEDOJ5 ( ICEDOJ5 )
 ,.ICEDOK3 ( ICEDOK3 ) ,.ICEDOL1 ( ICEDOL1 ) ,.ICEDOH8 ( ICEDOH8 ) ,.ICEDOJ4 ( ICEDOJ4 ) ,.ICEDOK2 ( ICEDOK2 ) ,.ICEDOL0 ( ICEDOL0 )
 ,.ICEDOJ31 ( ICEDOJ31 ) ,.ICEDOJ23 ( ICEDOJ23 ) ,.ICEDOJ15 ( ICEDOJ15 ) ,.ICEDOK11 ( ICEDOK11 ) ,.ICEDOJ30 ( ICEDOJ30 ) ,.ICEDOJ22 ( ICEDOJ22 )
 ,.ICEDOJ14 ( ICEDOJ14 ) ,.ICEDOK10 ( ICEDOK10 ) ,.ICEDOJ29 ( ICEDOJ29 ) ,.ICEDOK25 ( ICEDOK25 ) ,.ICEDOK17 ( ICEDOK17 ) ,.ICEDOL21 ( ICEDOL21 )
 ,.ICEDOL13 ( ICEDOL13 ) ,.ICEDOJ28 ( ICEDOJ28 ) ,.ICEDOK24 ( ICEDOK24 ) ,.ICEDOK16 ( ICEDOK16 ) ,.ICEDOL20 ( ICEDOL20 ) ,.ICEDOL12 ( ICEDOL12 )
 ,.ICEDOJ27 ( ICEDOJ27 ) ,.ICEDOJ19 ( ICEDOJ19 ) ,.ICEDOK31 ( ICEDOK31 ) ,.ICEDOK23 ( ICEDOK23 ) ,.ICEDOK15 ( ICEDOK15 ) ,.ICEDOL11 ( ICEDOL11 )
 ,.ICEDOJ26 ( ICEDOJ26 ) ,.ICEDOJ18 ( ICEDOJ18 ) ,.ICEDOK30 ( ICEDOK30 ) ,.ICEDOK22 ( ICEDOK22 ) ,.ICEDOK14 ( ICEDOK14 ) ,.ICEDOL10 ( ICEDOL10 )
 ,.ICEDOJ25 ( ICEDOJ25 ) ,.ICEDOJ17 ( ICEDOJ17 ) ,.ICEDOK21 ( ICEDOK21 ) ,.ICEDOK13 ( ICEDOK13 ) ,.ICEDOJ24 ( ICEDOJ24 ) ,.ICEDOJ16 ( ICEDOJ16 )
 ,.ICEDOK20 ( ICEDOK20 ) ,.ICEDOK12 ( ICEDOK12 ) ,.ICEDOJ9 ( ICEDOJ9 ) ,.ICEDOK7 ( ICEDOK7 ) ,.ICEDOL5 ( ICEDOL5 ) ,.ICEDOM3 ( ICEDOM3 )
 ,.ICEDON1 ( ICEDON1 ) ,.ICEDOJ8 ( ICEDOJ8 ) ,.ICEDOK6 ( ICEDOK6 ) ,.ICEDOL4 ( ICEDOL4 ) ,.ICEDOM2 ( ICEDOM2 ) ,.ICEDON0 ( ICEDON0 )
 ,.ICEDOJ7 ( ICEDOJ7 ) ,.ICEDOK5 ( ICEDOK5 ) ,.ICEDOL3 ( ICEDOL3 ) ,.ICEDOM1 ( ICEDOM1 ) ,.ICEDOJ6 ( ICEDOJ6 ) ,.ICEDOK4 ( ICEDOK4 )
 ,.ICEDOL2 ( ICEDOL2 ) ,.ICEDOM0 ( ICEDOM0 ) ,.ICEDOK29 ( ICEDOK29 ) ,.ICEDOL25 ( ICEDOL25 ) ,.ICEDOL17 ( ICEDOL17 ) ,.ICEDOM21 ( ICEDOM21 )
 ,.ICEDOM13 ( ICEDOM13 ) ,.ICEDOK28 ( ICEDOK28 ) ,.ICEDOL24 ( ICEDOL24 ) ,.ICEDOL16 ( ICEDOL16 ) ,.ICEDOM20 ( ICEDOM20 ) ,.ICEDOM12 ( ICEDOM12 )
 ,.ICEDOK27 ( ICEDOK27 ) ,.ICEDOK19 ( ICEDOK19 ) ,.ICEDOL31 ( ICEDOL31 ) ,.ICEDOL23 ( ICEDOL23 ) ,.ICEDOL15 ( ICEDOL15 ) ,.ICEDOM11 ( ICEDOM11 )
 ,.ICEDOK26 ( ICEDOK26 ) ,.ICEDOK18 ( ICEDOK18 ) ,.ICEDOL30 ( ICEDOL30 ) ,.ICEDOL22 ( ICEDOL22 ) ,.ICEDOL14 ( ICEDOL14 ) ,.ICEDOM10 ( ICEDOM10 )
 ,.ICEDOK9 ( ICEDOK9 ) ,.ICEDOL7 ( ICEDOL7 ) ,.ICEDOM5 ( ICEDOM5 ) ,.ICEDON3 ( ICEDON3 ) ,.ICEDOK8 ( ICEDOK8 ) ,.ICEDOL6 ( ICEDOL6 )
 ,.ICEDOM4 ( ICEDOM4 ) ,.ICEDON2 ( ICEDON2 ) ,.ICEDOL29 ( ICEDOL29 ) ,.ICEDOM25 ( ICEDOM25 ) ,.ICEDOM17 ( ICEDOM17 ) ,.ICEDON21 ( ICEDON21 )
 ,.ICEDON13 ( ICEDON13 ) ,.ICEDOL28 ( ICEDOL28 ) ,.ICEDOM24 ( ICEDOM24 ) ,.ICEDOM16 ( ICEDOM16 ) ,.ICEDON20 ( ICEDON20 ) ,.ICEDON12 ( ICEDON12 )
 ,.ICEDOL27 ( ICEDOL27 ) ,.ICEDOL19 ( ICEDOL19 ) ,.ICEDOM31 ( ICEDOM31 ) ,.ICEDOM23 ( ICEDOM23 ) ,.ICEDOM15 ( ICEDOM15 ) ,.ICEDON11 ( ICEDON11 )
 ,.ICEDOL26 ( ICEDOL26 ) ,.ICEDOL18 ( ICEDOL18 ) ,.ICEDOM30 ( ICEDOM30 ) ,.ICEDOM22 ( ICEDOM22 ) ,.ICEDOM14 ( ICEDOM14 ) ,.ICEDON10 ( ICEDON10 )
 ,.ICEDOL9 ( ICEDOL9 ) ,.ICEDOM7 ( ICEDOM7 ) ,.ICEDON5 ( ICEDON5 ) ,.ICEDOP1 ( ICEDOP1 ) ,.ICEDOL8 ( ICEDOL8 ) ,.ICEDOM6 ( ICEDOM6 )
 ,.ICEDON4 ( ICEDON4 ) ,.ICEDOP0 ( ICEDOP0 ) ,.ICEDOM29 ( ICEDOM29 ) ,.ICEDON25 ( ICEDON25 ) ,.ICEDON17 ( ICEDON17 ) ,.ICEDOM28 ( ICEDOM28 )
 ,.ICEDON24 ( ICEDON24 ) ,.ICEDON16 ( ICEDON16 ) ,.ICEDOM27 ( ICEDOM27 ) ,.ICEDOM19 ( ICEDOM19 ) ,.ICEDON31 ( ICEDON31 ) ,.ICEDON23 ( ICEDON23 )
 ,.ICEDON15 ( ICEDON15 ) ,.ICEDOM26 ( ICEDOM26 ) ,.ICEDOM18 ( ICEDOM18 ) ,.ICEDON30 ( ICEDON30 ) ,.ICEDON22 ( ICEDON22 ) ,.ICEDON14 ( ICEDON14 )
 ,.ICEDOM9 ( ICEDOM9 ) ,.ICEDON7 ( ICEDON7 ) ,.ICEDOP3 ( ICEDOP3 ) ,.ICEDOQ1 ( ICEDOQ1 ) ,.ICEDOM8 ( ICEDOM8 ) ,.ICEDON6 ( ICEDON6 )
 ,.ICEDOP2 ( ICEDOP2 ) ,.ICEDOQ0 ( ICEDOQ0 ) ,.ICEDON29 ( ICEDON29 ) ,.ICEDOP21 ( ICEDOP21 ) ,.ICEDOP13 ( ICEDOP13 ) ,.ICEDON28 ( ICEDON28 )
 ,.ICEDOP20 ( ICEDOP20 ) ,.ICEDOP12 ( ICEDOP12 ) ,.ICEDON27 ( ICEDON27 ) ,.ICEDON19 ( ICEDON19 ) ,.ICEDOP11 ( ICEDOP11 ) ,.ICEDON26 ( ICEDON26 )
 ,.ICEDON18 ( ICEDON18 ) ,.ICEDOP10 ( ICEDOP10 ) ,.ICEDON9 ( ICEDON9 ) ,.ICEDOP5 ( ICEDOP5 ) ,.ICEDOQ3 ( ICEDOQ3 ) ,.ICEDOR1 ( ICEDOR1 )
 ,.ICEDON8 ( ICEDON8 ) ,.ICEDOP4 ( ICEDOP4 ) ,.ICEDOQ2 ( ICEDOQ2 ) ,.ICEDOR0 ( ICEDOR0 ) ,.ICEDOP31 ( ICEDOP31 ) ,.ICEDOP23 ( ICEDOP23 )
 ,.ICEDOP15 ( ICEDOP15 ) ,.ICEDOQ11 ( ICEDOQ11 ) ,.ICEDOP30 ( ICEDOP30 ) ,.ICEDOP22 ( ICEDOP22 ) ,.ICEDOP14 ( ICEDOP14 ) ,.ICEDOQ10 ( ICEDOQ10 )
 ,.ICEDOP29 ( ICEDOP29 ) ,.ICEDOQ25 ( ICEDOQ25 ) ,.ICEDOQ17 ( ICEDOQ17 ) ,.ICEDOR21 ( ICEDOR21 ) ,.ICEDOR13 ( ICEDOR13 ) ,.ICEDOP28 ( ICEDOP28 )
 ,.ICEDOQ24 ( ICEDOQ24 ) ,.ICEDOQ16 ( ICEDOQ16 ) ,.ICEDOR20 ( ICEDOR20 ) ,.ICEDOR12 ( ICEDOR12 ) ,.ICEDOP27 ( ICEDOP27 ) ,.ICEDOP19 ( ICEDOP19 )
 ,.ICEDOQ31 ( ICEDOQ31 ) ,.ICEDOQ23 ( ICEDOQ23 ) ,.ICEDOQ15 ( ICEDOQ15 ) ,.ICEDOR11 ( ICEDOR11 ) ,.ICEDOP26 ( ICEDOP26 ) ,.ICEDOP18 ( ICEDOP18 )
 ,.ICEDOQ30 ( ICEDOQ30 ) ,.ICEDOQ22 ( ICEDOQ22 ) ,.ICEDOQ14 ( ICEDOQ14 ) ,.ICEDOR10 ( ICEDOR10 ) ,.ICEDOP25 ( ICEDOP25 ) ,.ICEDOP17 ( ICEDOP17 )
 ,.ICEDOQ21 ( ICEDOQ21 ) ,.ICEDOQ13 ( ICEDOQ13 ) ,.ICEDOP24 ( ICEDOP24 ) ,.ICEDOP16 ( ICEDOP16 ) ,.ICEDOQ20 ( ICEDOQ20 ) ,.ICEDOQ12 ( ICEDOQ12 )
 ,.ICEDOP9 ( ICEDOP9 ) ,.ICEDOQ7 ( ICEDOQ7 ) ,.ICEDOR5 ( ICEDOR5 ) ,.ICEDOS3 ( ICEDOS3 ) ,.ICEDOT1 ( ICEDOT1 ) ,.ICEDOP8 ( ICEDOP8 )
 ,.ICEDOQ6 ( ICEDOQ6 ) ,.ICEDOR4 ( ICEDOR4 ) ,.ICEDOS2 ( ICEDOS2 ) ,.ICEDOT0 ( ICEDOT0 ) ,.ICEDOP7 ( ICEDOP7 ) ,.ICEDOQ5 ( ICEDOQ5 )
 ,.ICEDOR3 ( ICEDOR3 ) ,.ICEDOS1 ( ICEDOS1 ) ,.ICEDOP6 ( ICEDOP6 ) ,.ICEDOQ4 ( ICEDOQ4 ) ,.ICEDOR2 ( ICEDOR2 ) ,.ICEDOS0 ( ICEDOS0 )
 ,.ICEDOQ29 ( ICEDOQ29 ) ,.ICEDOR25 ( ICEDOR25 ) ,.ICEDOR17 ( ICEDOR17 ) ,.ICEDOS21 ( ICEDOS21 ) ,.ICEDOS13 ( ICEDOS13 ) ,.ICEDOQ28 ( ICEDOQ28 )
 ,.ICEDOR24 ( ICEDOR24 ) ,.ICEDOR16 ( ICEDOR16 ) ,.ICEDOS20 ( ICEDOS20 ) ,.ICEDOS12 ( ICEDOS12 ) ,.ICEDOQ27 ( ICEDOQ27 ) ,.ICEDOQ19 ( ICEDOQ19 )
 ,.ICEDOR31 ( ICEDOR31 ) ,.ICEDOR23 ( ICEDOR23 ) ,.ICEDOR15 ( ICEDOR15 ) ,.ICEDOS11 ( ICEDOS11 ) ,.ICEDOQ26 ( ICEDOQ26 ) ,.ICEDOQ18 ( ICEDOQ18 )
 ,.ICEDOR30 ( ICEDOR30 ) ,.ICEDOR22 ( ICEDOR22 ) ,.ICEDOR14 ( ICEDOR14 ) ,.ICEDOS10 ( ICEDOS10 ) ,.ICEDOQ9 ( ICEDOQ9 ) ,.ICEDOR7 ( ICEDOR7 )
 ,.ICEDOS5 ( ICEDOS5 ) ,.ICEDOT3 ( ICEDOT3 ) ,.ICEDOU1 ( ICEDOU1 ) ,.ICEDOQ8 ( ICEDOQ8 ) ,.ICEDOR6 ( ICEDOR6 ) ,.ICEDOS4 ( ICEDOS4 )
 ,.ICEDOT2 ( ICEDOT2 ) ,.ICEDOU0 ( ICEDOU0 ) ,.ICEDOR29 ( ICEDOR29 ) ,.ICEDOS25 ( ICEDOS25 ) ,.ICEDOS17 ( ICEDOS17 ) ,.ICEDOT21 ( ICEDOT21 )
 ,.ICEDOT13 ( ICEDOT13 ) ,.ICEDOR28 ( ICEDOR28 ) ,.ICEDOS24 ( ICEDOS24 ) ,.ICEDOS16 ( ICEDOS16 ) ,.ICEDOT20 ( ICEDOT20 ) ,.ICEDOT12 ( ICEDOT12 )
 ,.ICEDOR27 ( ICEDOR27 ) ,.ICEDOR19 ( ICEDOR19 ) ,.ICEDOS31 ( ICEDOS31 ) ,.ICEDOS23 ( ICEDOS23 ) ,.ICEDOS15 ( ICEDOS15 ) ,.ICEDOT11 ( ICEDOT11 )
 ,.ICEDOR26 ( ICEDOR26 ) ,.ICEDOR18 ( ICEDOR18 ) ,.ICEDOS30 ( ICEDOS30 ) ,.ICEDOS22 ( ICEDOS22 ) ,.ICEDOS14 ( ICEDOS14 ) ,.ICEDOT10 ( ICEDOT10 )
 ,.ICEDOR9 ( ICEDOR9 ) ,.ICEDOS7 ( ICEDOS7 ) ,.ICEDOT5 ( ICEDOT5 ) ,.ICEDOU3 ( ICEDOU3 ) ,.ICEDOR8 ( ICEDOR8 ) ,.ICEDOS6 ( ICEDOS6 )
 ,.ICEDOT4 ( ICEDOT4 ) ,.ICEDOU2 ( ICEDOU2 ) ,.ICEDOS29 ( ICEDOS29 ) ,.ICEDOT25 ( ICEDOT25 ) ,.ICEDOT17 ( ICEDOT17 ) ,.ICEDOU21 ( ICEDOU21 )
 ,.ICEDOU13 ( ICEDOU13 ) ,.ICEDOS28 ( ICEDOS28 ) ,.ICEDOT24 ( ICEDOT24 ) ,.ICEDOT16 ( ICEDOT16 ) ,.ICEDOU20 ( ICEDOU20 ) ,.ICEDOU12 ( ICEDOU12 )
 ,.ICEDOS27 ( ICEDOS27 ) ,.ICEDOS19 ( ICEDOS19 ) ,.ICEDOT31 ( ICEDOT31 ) ,.ICEDOT23 ( ICEDOT23 ) ,.ICEDOT15 ( ICEDOT15 ) ,.ICEDOU11 ( ICEDOU11 )
 ,.ICEDOS26 ( ICEDOS26 ) ,.ICEDOS18 ( ICEDOS18 ) ,.ICEDOT30 ( ICEDOT30 ) ,.ICEDOT22 ( ICEDOT22 ) ,.ICEDOT14 ( ICEDOT14 ) ,.ICEDOU10 ( ICEDOU10 )
 ,.ICEDOS9 ( ICEDOS9 ) ,.ICEDOT7 ( ICEDOT7 ) ,.ICEDOU5 ( ICEDOU5 ) ,.ICEDOS8 ( ICEDOS8 ) ,.ICEDOT6 ( ICEDOT6 ) ,.ICEDOU4 ( ICEDOU4 )
 ,.ICEDOT29 ( ICEDOT29 ) ,.ICEDOU25 ( ICEDOU25 ) ,.ICEDOU17 ( ICEDOU17 ) ,.ICEDOT28 ( ICEDOT28 ) ,.ICEDOU24 ( ICEDOU24 ) ,.ICEDOU16 ( ICEDOU16 )
 ,.ICEDOT27 ( ICEDOT27 ) ,.ICEDOT19 ( ICEDOT19 ) ,.ICEDOU31 ( ICEDOU31 ) ,.ICEDOU23 ( ICEDOU23 ) ,.ICEDOU15 ( ICEDOU15 ) ,.ICEDOT26 ( ICEDOT26 )
 ,.ICEDOT18 ( ICEDOT18 ) ,.ICEDOU30 ( ICEDOU30 ) ,.ICEDOU22 ( ICEDOU22 ) ,.ICEDOU14 ( ICEDOU14 ) ,.ICEDOT9 ( ICEDOT9 ) ,.ICEDOU7 ( ICEDOU7 )
 ,.ICEDOT8 ( ICEDOT8 ) ,.ICEDOU6 ( ICEDOU6 ) ,.ICEDOU29 ( ICEDOU29 ) ,.ICEDOU28 ( ICEDOU28 ) ,.ICEDOU27 ( ICEDOU27 ) ,.ICEDOU19 ( ICEDOU19 )
 ,.ICEDOU26 ( ICEDOU26 ) ,.ICEDOU18 ( ICEDOU18 ) ,.ICEDOU9 ( ICEDOU9 ) ,.ICEDOU8 ( ICEDOU8 ) ,.ICEDI31 ( ICEDI31 ) ,.ICEDI23 ( ICEDI23 )
 ,.ICEDI15 ( ICEDI15 ) ,.ICEDI30 ( ICEDI30 ) ,.ICEDI22 ( ICEDI22 ) ,.ICEDI14 ( ICEDI14 ) ,.ICEDI29 ( ICEDI29 ) ,.ICEDI28 ( ICEDI28 )
 ,.ICEDI27 ( ICEDI27 ) ,.ICEDI19 ( ICEDI19 ) ,.ICEDI26 ( ICEDI26 ) ,.ICEDI18 ( ICEDI18 ) ,.ICEDI25 ( ICEDI25 ) ,.ICEDI17 ( ICEDI17 )
 ,.ICEDI24 ( ICEDI24 ) ,.ICEDI16 ( ICEDI16 ) ,.ICEDI21 ( ICEDI21 ) ,.ICEDI13 ( ICEDI13 ) ,.ICEDI20 ( ICEDI20 ) ,.ICEDI12 ( ICEDI12 )
 ,.ICEDI11 ( ICEDI11 ) ,.ICEDI10 ( ICEDI10 ) ,.ICEDI9 ( ICEDI9 ) ,.ICEDI8 ( ICEDI8 ) ,.ICEDI7 ( ICEDI7 ) ,.ICEDI6 ( ICEDI6 )
 ,.ICEDI5 ( ICEDI5 ) ,.ICEDI4 ( ICEDI4 ) ,.ICEDI3 ( ICEDI3 ) ,.ICEDI2 ( ICEDI2 ) ,.ICEDI1 ( ICEDI1 ) ,.ICEDI0 ( ICEDI0 )
 ,.ICERD ( ICERD ) ,.ICEWR ( ICEWR ) ,.ICEIFA_PRE31 ( ICEIFA_PRE31 ) ,.ICEIFA_PRE23 ( ICEIFA_PRE23 ) ,.ICEIFA_PRE15 ( ICEIFA_PRE15 ) ,.ICEIFA_PRE30 ( ICEIFA_PRE30 )
 ,.ICEIFA_PRE22 ( ICEIFA_PRE22 ) ,.ICEIFA_PRE14 ( ICEIFA_PRE14 ) ,.ICEIFA_PRE29 ( ICEIFA_PRE29 ) ,.ICEIFA_PRE28 ( ICEIFA_PRE28 ) ,.ICEIFA_PRE27 ( ICEIFA_PRE27 ) ,.ICEIFA_PRE19 ( ICEIFA_PRE19 )
 ,.ICEIFA_PRE26 ( ICEIFA_PRE26 ) ,.ICEIFA_PRE18 ( ICEIFA_PRE18 ) ,.ICEIFA_PRE25 ( ICEIFA_PRE25 ) ,.ICEIFA_PRE17 ( ICEIFA_PRE17 ) ,.ICEIFA_PRE24 ( ICEIFA_PRE24 ) ,.ICEIFA_PRE16 ( ICEIFA_PRE16 )
 ,.ICEIFA_PRE21 ( ICEIFA_PRE21 ) ,.ICEIFA_PRE13 ( ICEIFA_PRE13 ) ,.ICEIFA_PRE20 ( ICEIFA_PRE20 ) ,.ICEIFA_PRE12 ( ICEIFA_PRE12 ) ,.ICEIFA_PRE11 ( ICEIFA_PRE11 ) ,.ICEIFA_PRE10 ( ICEIFA_PRE10 )
 ,.ICEIFA_PRE9 ( ICEIFA_PRE9 ) ,.ICEIFA_PRE8 ( ICEIFA_PRE8 ) ,.ICEIFA_PRE7 ( ICEIFA_PRE7 ) ,.ICEIFA_PRE6 ( ICEIFA_PRE6 ) ,.ICEIFA_PRE5 ( ICEIFA_PRE5 ) ,.ICEIFA_PRE4 ( ICEIFA_PRE4 )
 ,.ICEIFA_PRE3 ( ICEIFA_PRE3 ) ,.ICEIFA_PRE2 ( ICEIFA_PRE2 ) ,.ICEIFA_PRE1 ( ICEIFA_PRE1 ) ,.ICEIFA_PRE0 ( ICEIFA_PRE0 ) ,.ICEDI_PRE31 ( ICEDI_PRE31 ) ,.ICEDI_PRE23 ( ICEDI_PRE23 )
 ,.ICEDI_PRE15 ( ICEDI_PRE15 ) ,.ICEDI_PRE30 ( ICEDI_PRE30 ) ,.ICEDI_PRE22 ( ICEDI_PRE22 ) ,.ICEDI_PRE14 ( ICEDI_PRE14 ) ,.ICEDI_PRE29 ( ICEDI_PRE29 ) ,.ICEDI_PRE28 ( ICEDI_PRE28 )
 ,.ICEDI_PRE27 ( ICEDI_PRE27 ) ,.ICEDI_PRE19 ( ICEDI_PRE19 ) ,.ICEDI_PRE26 ( ICEDI_PRE26 ) ,.ICEDI_PRE18 ( ICEDI_PRE18 ) ,.ICEDI_PRE25 ( ICEDI_PRE25 ) ,.ICEDI_PRE17 ( ICEDI_PRE17 )
 ,.ICEDI_PRE24 ( ICEDI_PRE24 ) ,.ICEDI_PRE16 ( ICEDI_PRE16 ) ,.ICEDI_PRE21 ( ICEDI_PRE21 ) ,.ICEDI_PRE13 ( ICEDI_PRE13 ) ,.ICEDI_PRE20 ( ICEDI_PRE20 ) ,.ICEDI_PRE12 ( ICEDI_PRE12 )
 ,.ICEDI_PRE11 ( ICEDI_PRE11 ) ,.ICEDI_PRE10 ( ICEDI_PRE10 ) ,.ICEDI_PRE9 ( ICEDI_PRE9 ) ,.ICEDI_PRE8 ( ICEDI_PRE8 ) ,.ICEDI_PRE7 ( ICEDI_PRE7 ) ,.ICEDI_PRE6 ( ICEDI_PRE6 )
 ,.ICEDI_PRE5 ( ICEDI_PRE5 ) ,.ICEDI_PRE4 ( ICEDI_PRE4 ) ,.ICEDI_PRE3 ( ICEDI_PRE3 ) ,.ICEDI_PRE2 ( ICEDI_PRE2 ) ,.ICEDI_PRE1 ( ICEDI_PRE1 ) ,.ICEDI_PRE0 ( ICEDI_PRE0 )
 ,.ICERD_PRE ( ICERD_PRE ) ,.ICEWR_PRE ( ICEWR_PRE ) ,.BASECK ( BASECK ) ,.SVMOD ( SVMOD ) ,.ALT1 ( ALT1 ) ,.SLMEM ( SLMEM )
 ,.MA15 ( MA15 ) ,.MA14 ( MA14 ) ,.MA13 ( MA13 ) ,.MA12 ( MA12 ) ,.MA11 ( MA11 ) ,.MA10 ( MA10 )
 ,.MA9 ( MA9 ) ,.MA8 ( MA8 ) ,.MA3 ( MA3 ) ,.MA2 ( MA2 ) ,.MA1 ( MA1 ) ,.MA0 ( MA0 )
 ,.MDW15 ( MDW15 ) ,.MDW14 ( MDW14 ) ,.MDW13 ( MDW13 ) ,.MDW12 ( MDW12 ) ,.MDW11 ( MDW11 ) ,.MDW10 ( MDW10 )
 ,.MDW9 ( MDW9 ) ,.MDW8 ( MDW8 ) ,.MDW7 ( MDW7 ) ,.MDW6 ( MDW6 ) ,.MDW5 ( MDW5 ) ,.MDW4 ( MDW4 )
 ,.MDW3 ( MDW3 ) ,.MDW2 ( MDW2 ) ,.MDW1 ( MDW1 ) ,.MDW0 ( MDW0 ) ,.CPUWR ( CPUWR ) ,.CPURD ( CPURD )
 ,.WDOP ( WDOP ) ,.VDDLEV7 ( VDDLEV7 ) ,.VDDLEV6 ( VDDLEV6 ) ,.VDDLEV5 ( VDDLEV5 ) ,.VDDLEV4 ( VDDLEV4 ) ,.VDDLEV3 ( VDDLEV3 )
 ,.VDDLEV2 ( VDDLEV2 ) ,.VDDLEV1 ( VDDLEV1 ) ,.VDDLEV0 ( VDDLEV0 ) ,.USBIFWR ( USBIFWR ) ,.ICECSGREGU ( ICECSGREGU ) ,.PC19 ( PC19 )
 ,.PC18 ( PC18 ) ,.PC17 ( PC17 ) ,.PC16 ( PC16 ) ,.PC15 ( PC15 ) ,.PC14 ( PC14 ) ,.PC13 ( PC13 )
 ,.PC12 ( PC12 ) ,.PC11 ( PC11 ) ,.PC10 ( PC10 ) ,.PC9 ( PC9 ) ,.PC8 ( PC8 ) ,.PC7 ( PC7 )
 ,.PC6 ( PC6 ) ,.PC5 ( PC5 ) ,.PC4 ( PC4 ) ,.PC3 ( PC3 ) ,.PC2 ( PC2 ) ,.PC1 ( PC1 )
 ,.PC0 ( PC0 )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/resetctl.v
  RESETCTL resetctl (
   .ICEIFA31 ( ICEIFA_PRE31 ) ,.ICEIFA23 ( ICEIFA_PRE23 ) ,.ICEIFA15 ( ICEIFA_PRE15 ) ,.ICEIFA30 ( ICEIFA_PRE30 ) ,.ICEIFA22 ( ICEIFA_PRE22 ) ,.ICEIFA14 ( ICEIFA_PRE14 ) ,.ICEIFA29 ( ICEIFA_PRE29 )
 ,.ICEIFA28 ( ICEIFA_PRE28 ) ,.ICEIFA27 ( ICEIFA_PRE27 ) ,.ICEIFA19 ( ICEIFA_PRE19 ) ,.ICEIFA26 ( ICEIFA_PRE26 ) ,.ICEIFA18 ( ICEIFA_PRE18 ) ,.ICEIFA25 ( ICEIFA_PRE25 )
 ,.ICEIFA17 ( ICEIFA_PRE17 ) ,.ICEIFA24 ( ICEIFA_PRE24 ) ,.ICEIFA16 ( ICEIFA_PRE16 ) ,.ICEIFA21 ( ICEIFA_PRE21 ) ,.ICEIFA13 ( ICEIFA_PRE13 ) ,.ICEIFA20 ( ICEIFA_PRE20 )
 ,.ICEIFA12 ( ICEIFA_PRE12 ) ,.ICEIFA11 ( ICEIFA_PRE11 ) ,.ICEIFA10 ( ICEIFA_PRE10 ) ,.ICEIFA9 ( ICEIFA_PRE9 ) ,.ICEIFA8 ( ICEIFA_PRE8 ) ,.ICEIFA7 ( ICEIFA_PRE7 )
 ,.ICEIFA6 ( ICEIFA_PRE6 ) ,.ICEIFA5 ( ICEIFA_PRE5 ) ,.ICEIFA4 ( ICEIFA_PRE4 ) ,.ICEIFA3 ( ICEIFA_PRE3 ) ,.ICEIFA2 ( ICEIFA_PRE2 ) ,.ICEDI0 ( ICEDI_PRE0 )
 ,.ICEWR ( ICEWR_PRE ) ,.CLK30MHZ ( CLK30MHZ_GB ) ,.ICESYSRES_B ( EICESYSRES_B ) ,.ICECPURES_B ( EICECPURES_B ) ,.ICEDO31 ( ICEDOB31 ) ,.ICEDO23 ( ICEDOB23 )
 ,.ICEDO15 ( ICEDOB15 ) ,.ICEDO30 ( ICEDOB30 ) ,.ICEDO22 ( ICEDOB22 ) ,.ICEDO14 ( ICEDOB14 ) ,.ICEDO29 ( ICEDOB29 ) ,.ICEDO28 ( ICEDOB28 )
 ,.ICEDO27 ( ICEDOB27 ) ,.ICEDO19 ( ICEDOB19 ) ,.ICEDO26 ( ICEDOB26 ) ,.ICEDO18 ( ICEDOB18 ) ,.ICEDO25 ( ICEDOB25 ) ,.ICEDO17 ( ICEDOB17 )
 ,.ICEDO24 ( ICEDOB24 ) ,.ICEDO16 ( ICEDOB16 ) ,.ICEDO21 ( ICEDOB21 ) ,.ICEDO13 ( ICEDOB13 ) ,.ICEDO20 ( ICEDOB20 ) ,.ICEDO12 ( ICEDOB12 )
 ,.ICEDO11 ( ICEDOB11 ) ,.ICEDO10 ( ICEDOB10 ) ,.ICEDO9 ( ICEDOB9 ) ,.ICEDO8 ( ICEDOB8 ) ,.ICEDO7 ( ICEDOB7 ) ,.ICEDO6 ( ICEDOB6 )
 ,.ICEDO5 ( ICEDOB5 ) ,.ICEDO4 ( ICEDOB4 ) ,.ICEDO3 ( ICEDOB3 ) ,.ICEDO2 ( ICEDOB2 ) ,.ICEDO1 ( ICEDOB1 ) ,.ICEDO0 ( ICEDOB0 )
 ,.CLK60MHZ ( CLK60MHZ ) ,.SVMODUSER ( SVMODUSER ) ,.PSEUDORES ( PSEUDORES ) ,.RESET_B ( RESET_B ) ,.ICEMSKPOC ( ICEMSKPOC ) ,.ICEMSKTRST ( ICEMSKTRST )
 ,.ICEMSKICE ( ICEMSKICE ) ,.ICEMSKTRSTFLG ( ICEMSKTRSTFLG ) ,.PONRESB ( PONRESB ) ,.ICERESB ( ICERESB ) ,.POCRESB ( POCRESB ) ,.TARRESB ( TARRESB )
 ,.TARRESB_NORM ( TARRESB_NORM ) ,.SYSRSOUTB ( SYSRSOUTB ) ,.BRKFAIL14 ( BRKFAIL14 )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/clockctl.v
  CLOCKCTL clockctl (
   .LOCKFAIL31 ( LOCK240FAIL ) ,.LOCKFAIL23 ( LOCKFAIL23 ) ,.LOCKFAIL15 ( LOCKFAIL15 ) ,.ICEDO31 ( ICEDOC31 ) ,.ICEDO23 ( ICEDOC23 ) ,.ICEDO15 ( ICEDOC15 ) ,.ICEDO30 ( ICEDOC30 )
 ,.ICEDO22 ( ICEDOC22 ) ,.ICEDO14 ( ICEDOC14 ) ,.ICEDO29 ( ICEDOC29 ) ,.ICEDO28 ( ICEDOC28 ) ,.ICEDO27 ( ICEDOC27 ) ,.ICEDO19 ( ICEDOC19 )
 ,.ICEDO26 ( ICEDOC26 ) ,.ICEDO18 ( ICEDOC18 ) ,.ICEDO25 ( ICEDOC25 ) ,.ICEDO17 ( ICEDOC17 ) ,.ICEDO24 ( ICEDOC24 ) ,.ICEDO16 ( ICEDOC16 )
 ,.ICEDO21 ( ICEDOC21 ) ,.ICEDO13 ( ICEDOC13 ) ,.ICEDO20 ( ICEDOC20 ) ,.ICEDO12 ( ICEDOC12 ) ,.ICEDO11 ( ICEDOC11 ) ,.ICEDO10 ( ICEDOC10 )
 ,.ICEDO9 ( ICEDOC9 ) ,.ICEDO8 ( ICEDOC8 ) ,.ICEDO7 ( ICEDOC7 ) ,.ICEDO6 ( ICEDOC6 ) ,.ICEDO5 ( ICEDOC5 ) ,.ICEDO4 ( ICEDOC4 )
 ,.ICEDO3 ( ICEDOC3 ) ,.ICEDO2 ( ICEDOC2 ) ,.ICEDO1 ( ICEDOC1 ) ,.ICEDO0 ( ICEDOC0 ) ,.SYSRSOUTB ( SYSRSOUTB ) ,.PONRESB ( PONRESB )
 ,.ICEIFA31 ( ICEIFA31 ) ,.ICEIFA23 ( ICEIFA23 ) ,.ICEIFA15 ( ICEIFA15 ) ,.ICEIFA30 ( ICEIFA30 ) ,.ICEIFA22 ( ICEIFA22 ) ,.ICEIFA14 ( ICEIFA14 )
 ,.ICEIFA29 ( ICEIFA29 ) ,.ICEIFA28 ( ICEIFA28 ) ,.ICEIFA27 ( ICEIFA27 ) ,.ICEIFA19 ( ICEIFA19 ) ,.ICEIFA26 ( ICEIFA26 ) ,.ICEIFA18 ( ICEIFA18 )
 ,.ICEIFA25 ( ICEIFA25 ) ,.ICEIFA17 ( ICEIFA17 ) ,.ICEIFA24 ( ICEIFA24 ) ,.ICEIFA16 ( ICEIFA16 ) ,.ICEIFA21 ( ICEIFA21 ) ,.ICEIFA13 ( ICEIFA13 )
 ,.ICEIFA20 ( ICEIFA20 ) ,.ICEIFA12 ( ICEIFA12 ) ,.ICEIFA11 ( ICEIFA11 ) ,.ICEIFA10 ( ICEIFA10 ) ,.ICEIFA9 ( ICEIFA9 ) ,.ICEIFA8 ( ICEIFA8 )
 ,.ICEIFA7 ( ICEIFA7 ) ,.ICEIFA6 ( ICEIFA6 ) ,.ICEIFA5 ( ICEIFA5 ) ,.ICEIFA4 ( ICEIFA4 ) ,.ICEIFA3 ( ICEIFA3 ) ,.ICEIFA2 ( ICEIFA2 )
 ,.ICEIFA1 ( ICEIFA1 ) ,.ICEIFA0 ( ICEIFA0 ) ,.ICEDI31 ( ICEDI31 ) ,.ICEDI23 ( ICEDI23 ) ,.ICEDI15 ( ICEDI15 ) ,.ICEDI30 ( ICEDI30 )
 ,.ICEDI22 ( ICEDI22 ) ,.ICEDI14 ( ICEDI14 ) ,.ICEDI29 ( ICEDI29 ) ,.ICEDI28 ( ICEDI28 ) ,.ICEDI27 ( ICEDI27 ) ,.ICEDI19 ( ICEDI19 )
 ,.ICEDI26 ( ICEDI26 ) ,.ICEDI18 ( ICEDI18 ) ,.ICEDI25 ( ICEDI25 ) ,.ICEDI17 ( ICEDI17 ) ,.ICEDI24 ( ICEDI24 ) ,.ICEDI16 ( ICEDI16 )
 ,.ICEDI21 ( ICEDI21 ) ,.ICEDI13 ( ICEDI13 ) ,.ICEDI20 ( ICEDI20 ) ,.ICEDI12 ( ICEDI12 ) ,.ICEDI11 ( ICEDI11 ) ,.ICEDI10 ( ICEDI10 )
 ,.ICEDI9 ( ICEDI9 ) ,.ICEDI8 ( ICEDI8 ) ,.ICEDI7 ( ICEDI7 ) ,.ICEDI6 ( ICEDI6 ) ,.ICEDI5 ( ICEDI5 ) ,.ICEDI4 ( ICEDI4 )
 ,.ICEDI3 ( ICEDI3 ) ,.ICEDI2 ( ICEDI2 ) ,.ICEDI1 ( ICEDI1 ) ,.ICEDI0 ( ICEDI0 ) ,.ICEWR ( ICEWR ) ,.CLK30MHZ ( CLK30MHZ )
 ,.CLK60MHZ ( CLK60MHZ ) ,.CPUTMCLK ( CPUTMCLK ) ,.EVAOSCMCLK ( EVAOSCMCLK ) ,.CPUTSCLK ( CPUTSCLK ) ,.CPURCLK1SEL ( CPURCLK1SEL ) ,.CPUPRCLK2 ( CPUPRCLK2 )
 ,.CPUPRCLK3 ( CPUPRCLK3 ) ,.EVAOSCRCLK1 ( EVAOSCRCLK1 ) ,.EVAOSCRCLK2 ( EVAOSCRCLK2 ) ,.EVAOSCRCLK3 ( EVAOSCRCLK3 ) ,.CPUMCLK ( CPUMCLK ) ,.CPUSCLK ( CPUSCLK )
 ,.CPURCLK1 ( CPURCLK1 ) ,.CPURCLK2 ( CPURCLK2 ) ,.CPURCLK3 ( CPURCLK3 ) ,.CLK60MHZLOCK ( CLK60MHZLOCK ) ,.LOCKFAIL30 ( LOCKFAIL30 ) ,.LOCKFAIL22 ( LOCKFAIL22 )
 ,.LOCKFAIL14 ( LOCKFAIL14 ) ,.LOCKFAIL29 ( LOCKFAIL29 ) ,.LOCKFAIL28 ( LOCKFAIL28 ) ,.LOCKFAIL27 ( LOCKFAIL27 ) ,.LOCKFAIL19 ( LOCKFAIL19 ) ,.LOCKFAIL26 ( LOCKFAIL26 )
 ,.LOCKFAIL18 ( LOCKFAIL18 ) ,.LOCKFAIL25 ( LOCKFAIL25 ) ,.LOCKFAIL17 ( LOCKFAIL17 ) ,.LOCKFAIL24 ( LOCKFAIL24 ) ,.LOCKFAIL16 ( LOCKFAIL16 ) ,.LOCKFAIL21 ( LOCKFAIL21 )
 ,.LOCKFAIL13 ( LOCKFAIL13 ) ,.LOCKFAIL20 ( LOCKFAIL20 ) ,.LOCKFAIL12 ( LOCKFAIL12 ) ,.LOCKFAIL11 ( LOCKFAIL11 ) ,.LOCKFAIL10 ( LOCKFAIL10 ) ,.LOCKFAIL9 ( LOCKFAIL9 )
 ,.LOCKFAIL8 ( LOCKFAIL8 ) ,.LOCKFAIL7 ( LOCKFAIL7 ) ,.LOCKFAIL6 ( LOCKFAIL6 ) ,.LOCKFAIL5 ( LOCKFAIL5 )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/break.v
  BREAK break (
   .CPURESETB ( CPURSOUTB ) ,.BRKFAIL14SOURCE ( BRKFAIL14 ) ,.BRKTMOT2 ( DOWN ) ,.BRKTMOT3 ( DOWN ) ,.BRKTMOT4 ( DOWN ) ,.BRKTMOV0 ( BRKTMOVR ) ,.BRKTMOT5 ( DOWN )
 ,.BRKTMOV1 ( BRKTMOVC0 ) ,.BRKTMOT6 ( DOWN ) ,.BRKTMOV2 ( BRKTMOVC1 ) ,.BRKTMOV3 ( BRKTMOVN0 ) ,.BRKTMOV4 ( BRKTMOVN1 ) ,.BRKTMOV5 ( DOWN )
 ,.BRKTMOV6 ( DOWN ) ,.ICEDO31 ( ICEDOF31 ) ,.ICEDO23 ( ICEDOF23 ) ,.ICEDO15 ( ICEDOF15 ) ,.ICEDO30 ( ICEDOF30 ) ,.ICEDO22 ( ICEDOF22 )
 ,.ICEDO14 ( ICEDOF14 ) ,.ICEDO29 ( ICEDOF29 ) ,.ICEDO28 ( ICEDOF28 ) ,.ICEDO27 ( ICEDOF27 ) ,.ICEDO19 ( ICEDOF19 ) ,.ICEDO26 ( ICEDOF26 )
 ,.ICEDO18 ( ICEDOF18 ) ,.ICEDO25 ( ICEDOF25 ) ,.ICEDO17 ( ICEDOF17 ) ,.ICEDO24 ( ICEDOF24 ) ,.ICEDO16 ( ICEDOF16 ) ,.ICEDO21 ( ICEDOF21 )
 ,.ICEDO13 ( ICEDOF13 ) ,.ICEDO20 ( ICEDOF20 ) ,.ICEDO12 ( ICEDOF12 ) ,.ICEDO11 ( ICEDOF11 ) ,.ICEDO10 ( ICEDOF10 ) ,.ICEDO9 ( ICEDOF9 )
 ,.ICEDO8 ( ICEDOF8 ) ,.ICEDO7 ( ICEDOF7 ) ,.ICEDO6 ( ICEDOF6 ) ,.ICEDO5 ( ICEDOF5 ) ,.ICEDO4 ( ICEDOF4 ) ,.ICEDO3 ( ICEDOF3 )
 ,.ICEDO2 ( ICEDOF2 ) ,.ICEDO1 ( ICEDOF1 ) ,.ICEDO0 ( ICEDOF0 ) ,.ES3 ( EXMA3 ) ,.MA7 ( MA7 ) ,.ES2 ( EXMA2 )
 ,.MA6 ( MA6 ) ,.ES1 ( EXMA1 ) ,.MA5 ( MA5 ) ,.ES0 ( EXMA0 ) ,.MA4 ( MA4 ) ,.MDR15 ( BRKMDR15 )
 ,.MDR14 ( BRKMDR14 ) ,.MDR13 ( BRKMDR13 ) ,.MDR12 ( BRKMDR12 ) ,.MDR11 ( BRKMDR11 ) ,.MDR10 ( BRKMDR10 ) ,.MDR9 ( BRKMDR9 )
 ,.MDR8 ( BRKMDR8 ) ,.MDR7 ( BRKMDR7 ) ,.MDR6 ( BRKMDR6 ) ,.MDR5 ( BRKMDR5 ) ,.MDR4 ( BRKMDR4 ) ,.MDR3 ( BRKMDR3 )
 ,.MDR2 ( BRKMDR2 ) ,.MDR1 ( BRKMDR1 ) ,.MDR0 ( BRKMDR0 ) ,.SYSRSOUTB ( SYSRSOUTB ) ,.CLK60MHZ ( CLK60MHZ ) ,.ICEIFA31 ( ICEIFA31 )
 ,.ICEIFA23 ( ICEIFA23 ) ,.ICEIFA15 ( ICEIFA15 ) ,.ICEIFA30 ( ICEIFA30 ) ,.ICEIFA22 ( ICEIFA22 ) ,.ICEIFA14 ( ICEIFA14 ) ,.ICEIFA29 ( ICEIFA29 )
 ,.ICEIFA28 ( ICEIFA28 ) ,.ICEIFA27 ( ICEIFA27 ) ,.ICEIFA19 ( ICEIFA19 ) ,.ICEIFA26 ( ICEIFA26 ) ,.ICEIFA18 ( ICEIFA18 ) ,.ICEIFA25 ( ICEIFA25 )
 ,.ICEIFA17 ( ICEIFA17 ) ,.ICEIFA24 ( ICEIFA24 ) ,.ICEIFA16 ( ICEIFA16 ) ,.ICEIFA21 ( ICEIFA21 ) ,.ICEIFA13 ( ICEIFA13 ) ,.ICEIFA20 ( ICEIFA20 )
 ,.ICEIFA12 ( ICEIFA12 ) ,.ICEIFA11 ( ICEIFA11 ) ,.ICEIFA10 ( ICEIFA10 ) ,.ICEIFA9 ( ICEIFA9 ) ,.ICEIFA8 ( ICEIFA8 ) ,.ICEIFA7 ( ICEIFA7 )
 ,.ICEIFA6 ( ICEIFA6 ) ,.ICEIFA5 ( ICEIFA5 ) ,.ICEIFA4 ( ICEIFA4 ) ,.ICEIFA3 ( ICEIFA3 ) ,.ICEIFA2 ( ICEIFA2 ) ,.ICEIFA1 ( ICEIFA1 )
 ,.ICEIFA0 ( ICEIFA0 ) ,.ICEDI31 ( ICEDI31 ) ,.ICEDI23 ( ICEDI23 ) ,.ICEDI15 ( ICEDI15 ) ,.IDADR11 ( IDADR11 ) ,.ICEDI30 ( ICEDI30 )
 ,.ICEDI22 ( ICEDI22 ) ,.ICEDI14 ( ICEDI14 ) ,.IDADR10 ( IDADR10 ) ,.ICEDI29 ( ICEDI29 ) ,.ICEDI28 ( ICEDI28 ) ,.ICEDI27 ( ICEDI27 )
 ,.ICEDI19 ( ICEDI19 ) ,.IDADR15 ( IDADR15 ) ,.ICEDI26 ( ICEDI26 ) ,.ICEDI18 ( ICEDI18 ) ,.IDADR14 ( IDADR14 ) ,.ICEDI25 ( ICEDI25 )
 ,.ICEDI17 ( ICEDI17 ) ,.IDADR13 ( IDADR13 ) ,.ICEDI24 ( ICEDI24 ) ,.ICEDI16 ( ICEDI16 ) ,.IDADR12 ( IDADR12 ) ,.ICEDI21 ( ICEDI21 )
 ,.ICEDI13 ( ICEDI13 ) ,.ICEDI20 ( ICEDI20 ) ,.ICEDI12 ( ICEDI12 ) ,.ICEDI11 ( ICEDI11 ) ,.ICEDI10 ( ICEDI10 ) ,.ICEDI9 ( ICEDI9 )
 ,.IDADR7 ( IDADR7 ) ,.ICEDI8 ( ICEDI8 ) ,.IDADR6 ( IDADR6 ) ,.ICEDI7 ( ICEDI7 ) ,.IDADR5 ( IDADR5 ) ,.ICEDI6 ( ICEDI6 )
 ,.IDADR4 ( IDADR4 ) ,.ICEDI5 ( ICEDI5 ) ,.IDADR3 ( IDADR3 ) ,.ICEDI4 ( ICEDI4 ) ,.IDADR2 ( IDADR2 ) ,.ICEDI3 ( ICEDI3 )
 ,.IDADR1 ( IDADR1 ) ,.ICEDI2 ( ICEDI2 ) ,.IDADR0 ( IDADR0 ) ,.ICEDI1 ( ICEDI1 ) ,.ICEDI0 ( ICEDI0 ) ,.ICEWR ( ICEWR )
 ,.BASECK ( BASECK ) ,.SLMEM ( SLMEM ) ,.MA15 ( MA15 ) ,.MA14 ( MA14 ) ,.MA13 ( MA13 ) ,.MA12 ( MA12 )
 ,.MA11 ( MA11 ) ,.MA10 ( MA10 ) ,.MA9 ( MA9 ) ,.MA8 ( MA8 ) ,.MA3 ( MA3 ) ,.MA2 ( MA2 )
 ,.MA1 ( MA1 ) ,.MA0 ( MA0 ) ,.MDW15 ( MDW15 ) ,.MDW14 ( MDW14 ) ,.MDW13 ( MDW13 ) ,.MDW12 ( MDW12 )
 ,.MDW11 ( MDW11 ) ,.MDW10 ( MDW10 ) ,.MDW9 ( MDW9 ) ,.MDW8 ( MDW8 ) ,.MDW7 ( MDW7 ) ,.MDW6 ( MDW6 )
 ,.MDW5 ( MDW5 ) ,.MDW4 ( MDW4 ) ,.MDW3 ( MDW3 ) ,.MDW2 ( MDW2 ) ,.MDW1 ( MDW1 ) ,.MDW0 ( MDW0 )
 ,.CPUWR ( CPUWR ) ,.CPURD ( CPURD ) ,.SVMOD ( SVMOD ) ,.SVMODF ( SVMODF ) ,.HLTST ( HLTST ) ,.STPST ( STPST )
 ,.ALT1 ( ALT1 ) ,.SELFMODEDBG ( SELFMODEDBG ) ,.BRKFAIL0 ( BRKFAIL0 ) ,.BRKFAIL1 ( BRKFAIL1 ) ,.BRKFAIL2 ( BRKFAIL2 ) ,.BRKFAIL3 ( BRKFAIL3 )
 ,.BRKFAIL4 ( BRKFAIL4 ) ,.BRKFAIL5 ( BRKFAIL5 ) ,.BRKFAIL6 ( BRKFAIL6 ) ,.BRKFAIL7 ( BRKFAIL7 ) ,.BRKFAIL8 ( BRKFAIL8 ) ,.BRKFAIL9 ( BRKFAIL9 )
 ,.BRKFAIL10 ( BRKFAIL10 ) ,.BRKFAIL11 ( BRKFAIL11 ) ,.BRKFAIL12 ( BRKFAIL12 ) ,.BRKFAIL13 ( BRKFAIL13 ) ,.BRKFAIL15 ( BRKFAIL15 ) ,.SOFTBRK ( SOFTBRK )
 ,.BRKEDMM0 ( BRKEDMM0 ) ,.BRKEDMM1 ( BRKEDMM1 ) ,.BRKEDMM2 ( BRKEDMM2 ) ,.BRKEDMM3 ( BRKEDMM3 ) ,.BRKSNAP0 ( BRKSNAP0 ) ,.BRKSNAP1 ( BRKSNAP1 )
 ,.BRKSNAP2 ( BRKSNAP2 ) ,.BRKEVTF0 ( BRKEVTF0 ) ,.BRKEVTF1 ( BRKEVTF1 ) ,.BRKEVTF2 ( BRKEVTF2 ) ,.BRKEVTF3 ( BRKEVTF3 ) ,.BRKEVTF4 ( BRKEVTF4 )
 ,.BRKEVTF5 ( BRKEVTF5 ) ,.BRKEVTF6 ( BRKEVTF6 ) ,.BRKEVTF7 ( BRKEVTF7 ) ,.BRKEVTA0 ( BRKEVTA0 ) ,.BRKEVTA1 ( BRKEVTA1 ) ,.BRKEVTA2 ( BRKEVTA2 )
 ,.BRKEVTA3 ( BRKEVTA3 ) ,.BRKEVTA4 ( BRKEVTA4 ) ,.BRKEVTA5 ( BRKEVTA5 ) ,.BRKEVTA6 ( BRKEVTA6 ) ,.BRKEVTA7 ( BRKEVTA7 ) ,.BRKEVTL0 ( BRKEVTL0 )
 ,.BRKEVTL1 ( BRKEVTL1 ) ,.BRKTMOT0 ( BRKTMOT0 ) ,.BRKTMOT1 ( BRKTMOT1 ) ,.BRKTRAFL ( BRKTRAFL ) ,.BRKTRADY ( BRKTRADY ) ,.STBRELESV ( STBRELESV )
 ,.SVI ( SVI ) ,.SVVCOUT7 ( SVVCOUT7 ) ,.SVVCOUT6 ( SVVCOUT6 ) ,.SVVCOUT5 ( SVVCOUT5 ) ,.SVVCOUT4 ( SVVCOUT4 ) ,.SVVCOUT3 ( SVVCOUT3 )
 ,.SVVCOUT2 ( SVVCOUT2 ) ,.SVVCOUT1 ( SVVCOUT1 ) ,.SVVCOUT0 ( SVVCOUT0 ) ,.SVINTACK ( SVINTACK ) ,.PCWAITF ( PCWAITF ) ,.SVMODI ( SVMODI )
 ,.SVMODUSER ( SVMODUSER ) ,.SVMODOPBRK ( SVMODOPBRK ) ,.SVMODIPERI1 ( SVMODIPERI1 ) ,.SVMODIPERI2 ( SVMODIPERI2 ) ,.STEP ( STEP ) ,.IDADR9 ( IDADR9 )
 ,.IDADR8 ( IDADR8 )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/tracev1.v
  TRACE trace (
   .CLK30MHZ ( CLK30MHZ_GB ) ,.ICEDO31 ( ICEDOG31 ) ,.ICEDO23 ( ICEDOG23 ) ,.ICEDO15 ( ICEDOG15 ) ,.ICEDO30 ( ICEDOG30 ) ,.ICEDO22 ( ICEDOG22 ) ,.ICEDO14 ( ICEDOG14 )
 ,.ICEDO29 ( ICEDOG29 ) ,.ICEDO28 ( ICEDOG28 ) ,.ICEDO27 ( ICEDOG27 ) ,.ICEDO19 ( ICEDOG19 ) ,.ICEDO26 ( ICEDOG26 ) ,.ICEDO18 ( ICEDOG18 )
 ,.ICEDO25 ( ICEDOG25 ) ,.ICEDO17 ( ICEDOG17 ) ,.ICEDO24 ( ICEDOG24 ) ,.ICEDO16 ( ICEDOG16 ) ,.ICEDO21 ( ICEDOG21 ) ,.ICEDO13 ( ICEDOG13 )
 ,.ICEDO20 ( ICEDOG20 ) ,.ICEDO12 ( ICEDOG12 ) ,.ICEDO11 ( ICEDOG11 ) ,.ICEDO10 ( ICEDOG10 ) ,.ICEDO9 ( ICEDOG9 ) ,.ICEDO8 ( ICEDOG8 )
 ,.ICEDO7 ( ICEDOG7 ) ,.ICEDO6 ( ICEDOG6 ) ,.ICEDO5 ( ICEDOG5 ) ,.ICEDO4 ( ICEDOG4 ) ,.ICEDO3 ( ICEDOG3 ) ,.ICEDO2 ( ICEDOG2 )
 ,.ICEDO1 ( ICEDOG1 ) ,.ICEDO0 ( ICEDOG0 ) ,.ICEIFA31 ( ICEIFA31 ) ,.ICEIFA23 ( ICEIFA23 ) ,.ICEIFA15 ( ICEIFA15 ) ,.ICEIFA30 ( ICEIFA30 )
 ,.ICEIFA22 ( ICEIFA22 ) ,.ICEIFA14 ( ICEIFA14 ) ,.ICEIFA29 ( ICEIFA29 ) ,.ICEIFA28 ( ICEIFA28 ) ,.ICEIFA27 ( ICEIFA27 ) ,.ICEIFA19 ( ICEIFA19 )
 ,.ICEIFA26 ( ICEIFA26 ) ,.ICEIFA18 ( ICEIFA18 ) ,.ICEIFA25 ( ICEIFA25 ) ,.ICEIFA17 ( ICEIFA17 ) ,.ICEIFA24 ( ICEIFA24 ) ,.ICEIFA16 ( ICEIFA16 )
 ,.ICEIFA21 ( ICEIFA21 ) ,.ICEIFA13 ( ICEIFA13 ) ,.ICEIFA20 ( ICEIFA20 ) ,.ICEIFA12 ( ICEIFA12 ) ,.ICEIFA11 ( ICEIFA11 ) ,.ICEIFA10 ( ICEIFA10 )
 ,.ICEIFA9 ( ICEIFA9 ) ,.ICEIFA8 ( ICEIFA8 ) ,.ICEIFA7 ( ICEIFA7 ) ,.ICEIFA6 ( ICEIFA6 ) ,.ICEIFA5 ( ICEIFA5 ) ,.ICEIFA4 ( ICEIFA4 )
 ,.ICEIFA3 ( ICEIFA3 ) ,.ICEIFA2 ( ICEIFA2 ) ,.ICEDI31 ( ICEDI31 ) ,.ICEDI23 ( ICEDI23 ) ,.ICEDI15 ( ICEDI15 ) ,.IDADR11 ( IDADR11 )
 ,.ICEDI30 ( ICEDI30 ) ,.ICEDI22 ( ICEDI22 ) ,.ICEDI14 ( ICEDI14 ) ,.IDADR10 ( IDADR10 ) ,.ICEDI29 ( ICEDI29 ) ,.IDADR25 ( IDADR25 )
 ,.IDADR17 ( IDADR17 ) ,.ICEDI28 ( ICEDI28 ) ,.IDADR24 ( IDADR24 ) ,.IDADR16 ( IDADR16 ) ,.ICEDI27 ( ICEDI27 ) ,.ICEDI19 ( ICEDI19 )
 ,.IDADR31 ( IDADR31 ) ,.IDADR23 ( IDADR23 ) ,.IDADR15 ( IDADR15 ) ,.ICEDI26 ( ICEDI26 ) ,.ICEDI18 ( ICEDI18 ) ,.IDADR30 ( IDADR30 )
 ,.IDADR22 ( IDADR22 ) ,.IDADR14 ( IDADR14 ) ,.ICEDI25 ( ICEDI25 ) ,.ICEDI17 ( ICEDI17 ) ,.IDADR21 ( IDADR21 ) ,.IDADR13 ( IDADR13 )
 ,.ICEDI24 ( ICEDI24 ) ,.ICEDI16 ( ICEDI16 ) ,.IDADR20 ( IDADR20 ) ,.IDADR12 ( IDADR12 ) ,.ICEDI21 ( ICEDI21 ) ,.ICEDI13 ( ICEDI13 )
 ,.ICEDI20 ( ICEDI20 ) ,.ICEDI12 ( ICEDI12 ) ,.ICEDI11 ( ICEDI11 ) ,.ICEDI10 ( ICEDI10 ) ,.ICEDI9 ( ICEDI9 ) ,.IDADR7 ( IDADR7 )
 ,.ICEDI8 ( ICEDI8 ) ,.IDADR6 ( IDADR6 ) ,.ICEDI7 ( ICEDI7 ) ,.IDADR5 ( IDADR5 ) ,.ICEDI6 ( ICEDI6 ) ,.IDADR4 ( IDADR4 )
 ,.ICEDI5 ( ICEDI5 ) ,.IDADR3 ( IDADR3 ) ,.ICEDI4 ( ICEDI4 ) ,.IDADR2 ( IDADR2 ) ,.ICEDI3 ( ICEDI3 ) ,.IDADR1 ( IDADR1 )
 ,.ICEDI2 ( ICEDI2 ) ,.IDADR0 ( IDADR0 ) ,.ICEDI1 ( ICEDI1 ) ,.ICEDI0 ( ICEDI0 ) ,.ICEWR ( ICEWR ) ,.PC19 ( PC19 )
 ,.PC18 ( PC18 ) ,.PC17 ( PC17 ) ,.PC16 ( PC16 ) ,.PC15 ( PC15 ) ,.PC14 ( PC14 ) ,.PC13 ( PC13 )
 ,.PC12 ( PC12 ) ,.PC11 ( PC11 ) ,.PC10 ( PC10 ) ,.PC9 ( PC9 ) ,.PC8 ( PC8 ) ,.PC7 ( PC7 )
 ,.PC6 ( PC6 ) ,.PC5 ( PC5 ) ,.PC4 ( PC4 ) ,.PC3 ( PC3 ) ,.PC2 ( PC2 ) ,.PC1 ( PC1 )
 ,.PC0 ( PC0 ) ,.IDADR29 ( IDADR29 ) ,.IDADR28 ( IDADR28 ) ,.IDADR27 ( IDADR27 ) ,.IDADR19 ( IDADR19 ) ,.IDADR26 ( IDADR26 )
 ,.IDADR18 ( IDADR18 ) ,.IDADR9 ( IDADR9 ) ,.IDADR8 ( IDADR8 ) ,.STAGEADR1 ( STAGEADR1 ) ,.STAGEADR0 ( STAGEADR0 ) ,.PREFIX ( PREFIX )
 ,.FLREAD ( FLREAD ) ,.IMDR10 ( IMDR10 ) ,.FLREADB3 ( FLREADB3 ) ,.FLREADB2 ( FLREADB2 ) ,.FLREADB1 ( FLREADB1 ) ,.FLREADB0 ( FLREADB0 )
 ,.EROMPD31 ( EROMPD31 ) ,.EROMPD23 ( EROMPD23 ) ,.EROMPD15 ( EROMPD15 ) ,.EROMPD30 ( EROMPD30 ) ,.EROMPD22 ( EROMPD22 ) ,.EROMPD14 ( EROMPD14 )
 ,.EROMPD29 ( EROMPD29 ) ,.EROMPD28 ( EROMPD28 ) ,.EROMPD27 ( EROMPD27 ) ,.EROMPD19 ( EROMPD19 ) ,.EROMPD26 ( EROMPD26 ) ,.EROMPD18 ( EROMPD18 )
 ,.EROMPD25 ( EROMPD25 ) ,.EROMPD17 ( EROMPD17 ) ,.EROMPD24 ( EROMPD24 ) ,.EROMPD16 ( EROMPD16 ) ,.EROMPD21 ( EROMPD21 ) ,.EROMPD13 ( EROMPD13 )
 ,.EROMPD20 ( EROMPD20 ) ,.EROMPD12 ( EROMPD12 ) ,.EROMPD11 ( EROMPD11 ) ,.EROMPD10 ( EROMPD10 ) ,.EROMPD9 ( EROMPD9 ) ,.EROMPD8 ( EROMPD8 )
 ,.EROMPD7 ( EROMPD7 ) ,.EROMPD6 ( EROMPD6 ) ,.EROMPD5 ( EROMPD5 ) ,.EROMPD4 ( EROMPD4 ) ,.EROMPD3 ( EROMPD3 ) ,.EROMPD2 ( EROMPD2 )
 ,.EROMPD1 ( EROMPD1 ) ,.EROMPD0 ( EROMPD0 ) ,.PCWAITF ( PCWAITF ) ,.WAITEXM ( WAITEXM ) ,.OCDWAIT ( OCDWAIT ) ,.SKIPEXE ( SKIPEXE )
 ,.FCHRAM ( FCHRAM ) ,.CPUMASK ( CPUMASK ) ,.EXMA3 ( EXMA3 ) ,.TAG21 ( TAG21 ) ,.TAG13 ( TAG13 ) ,.EXMA2 ( EXMA2 )
 ,.TAG20 ( TAG20 ) ,.TAG12 ( TAG12 ) ,.EXMA1 ( EXMA1 ) ,.TAG11 ( TAG11 ) ,.EXMA0 ( EXMA0 ) ,.TAG10 ( TAG10 )
 ,.MA15 ( MA15 ) ,.MA14 ( MA14 ) ,.MA13 ( MA13 ) ,.MA12 ( MA12 ) ,.MA11 ( MA11 ) ,.MA10 ( MA10 )
 ,.MA9 ( MA9 ) ,.MA8 ( MA8 ) ,.MA7 ( MA7 ) ,.MA6 ( MA6 ) ,.MA5 ( MA5 ) ,.MA4 ( MA4 )
 ,.MA3 ( MA3 ) ,.MA2 ( MA2 ) ,.MA1 ( MA1 ) ,.MA0 ( MA0 ) ,.IMDR15 ( IMDR15 ) ,.IMDR14 ( IMDR14 )
 ,.IMDR13 ( IMDR13 ) ,.IMDR12 ( IMDR12 ) ,.IMDR11 ( IMDR11 ) ,.IMDR9 ( IMDR9 ) ,.IMDR8 ( IMDR8 ) ,.IMDR7 ( IMDR7 )
 ,.MDW15 ( MDW15 ) ,.IMDR6 ( IMDR6 ) ,.MDW14 ( MDW14 ) ,.IMDR5 ( IMDR5 ) ,.MDW13 ( MDW13 ) ,.IMDR4 ( IMDR4 )
 ,.MDW12 ( MDW12 ) ,.IMDR3 ( IMDR3 ) ,.MDW11 ( MDW11 ) ,.IMDR2 ( IMDR2 ) ,.MDW10 ( MDW10 ) ,.IMDR1 ( IMDR1 )
 ,.IMDR0 ( IMDR0 ) ,.TRACEMDR15 ( TRACEMDR15 ) ,.TRACEMDR14 ( TRACEMDR14 ) ,.TRACEMDR13 ( TRACEMDR13 ) ,.TRACEMDR12 ( TRACEMDR12 ) ,.TRACEMDR11 ( TRACEMDR11 )
 ,.TRACEMDR10 ( TRACEMDR10 ) ,.TRACEMDR9 ( TRACEMDR9 ) ,.TRACEMDR8 ( TRACEMDR8 ) ,.TRACEMDR7 ( TRACEMDR7 ) ,.TRACEMDR6 ( TRACEMDR6 ) ,.TRACEMDR5 ( TRACEMDR5 )
 ,.TRACEMDR4 ( TRACEMDR4 ) ,.TRACEMDR3 ( TRACEMDR3 ) ,.TRACEMDR2 ( TRACEMDR2 ) ,.TRACEMDR1 ( TRACEMDR1 ) ,.TRACEMDR0 ( TRACEMDR0 ) ,.MDW9 ( MDW9 )
 ,.MDW8 ( MDW8 ) ,.MDW7 ( MDW7 ) ,.MDW6 ( MDW6 ) ,.MDW5 ( MDW5 ) ,.MDW4 ( MDW4 ) ,.MDW3 ( MDW3 )
 ,.MDW2 ( MDW2 ) ,.MDW1 ( MDW1 ) ,.MDW0 ( MDW0 ) ,.CPURD ( CPURD ) ,.CPUWR ( CPUWR ) ,.WDOP ( WDOP )
 ,.BASECK ( BASECK ) ,.ALT1 ( ALT1 ) ,.SVMOD ( SVMOD ) ,.SVMODUSER ( SVMODUSER ) ,.SELFMODE ( SELFMODE ) ,.SELFMODEDBG ( SELFMODEDBG )
 ,.SELEXMPC ( SELEXMPC ) ,.SELRAMPC ( SELRAMPC ) ,.SELROMPC ( SELROMPC ) ,.SELBRAMPC ( SELBRAMPC ) ,.SELBFAPC ( SELBFAPC ) ,.TAG31 ( TAG31 )
 ,.TAG23 ( TAG23 ) ,.TAG15 ( TAG15 ) ,.TAG30 ( TAG30 ) ,.TAG22 ( TAG22 ) ,.TAG14 ( TAG14 ) ,.TAG29 ( TAG29 )
 ,.TAG28 ( TAG28 ) ,.TAG27 ( TAG27 ) ,.TAG19 ( TAG19 ) ,.TAG26 ( TAG26 ) ,.TAG18 ( TAG18 ) ,.TAG25 ( TAG25 )
 ,.TAG17 ( TAG17 ) ,.TAG24 ( TAG24 ) ,.TAG16 ( TAG16 ) ,.TAG9 ( TAG9 ) ,.TAG8 ( TAG8 ) ,.TAG7 ( TAG7 )
 ,.TAG6 ( TAG6 ) ,.TAG5 ( TAG5 ) ,.TAG4 ( TAG4 ) ,.TAG3 ( TAG3 ) ,.TAG2 ( TAG2 ) ,.TAG1 ( TAG1 )
 ,.TAG0 ( TAG0 ) ,.TAGOVF ( TAGOVF ) ,.CLK60MHZ ( CLK60MHZ ) ,.SYSRSOUTB ( SYSRSOUTB ) ,.ICERESB ( ICERESB ) ,.CPURSOUTB ( CPURSOUTB )
 ,.TARRESB_NORM ( TARRESB_NORM ) ,.ICEMSKICE ( ICEMSKICE ) ,.ICEMSKTRST ( ICEMSKTRST ) ,.STEP ( STEP ) ,.INTACK ( INTACK ) ,.DMAACK ( DMAACK )
 ,.BRKTRADY ( BRKTRADY ) ,.BRKTRAFL ( BRKTRAFL ) ,.EVD01 ( EVD01 ) ,.EVD02 ( EVD02 ) ,.EVD10 ( EVD10 ) ,.EVD03 ( EVD03 )
 ,.EVD04 ( EVD04 ) ,.EVD05 ( EVD05 ) ,.EVD06 ( EVD06 ) ,.EVD07 ( EVD07 ) ,.EVD08 ( EVD08 ) ,.EVD09 ( EVD09 )
 ,.TRCON ( TRCON ) ,.MONITRC ( MONITRC ) ,.TRCMD ( TRCMD ) ,.TMEMWAIT ( TMEMWAIT ) ,.TMEMA16 ( TMEMA16 ) ,.TMEMA15 ( TMEMA15 )
 ,.TMEMA14 ( TMEMA14 ) ,.TMEMA13 ( TMEMA13 ) ,.TMEMA12 ( TMEMA12 ) ,.TMEMA11 ( TMEMA11 ) ,.TMEMA10 ( TMEMA10 ) ,.TMEMA9 ( TMEMA9 )
 ,.TMEMD3 ( TMEMD3 ) ,.TMEMA8 ( TMEMA8 ) ,.TMEMD2 ( TMEMD2 ) ,.TMEMA7 ( TMEMA7 ) ,.TMEMD1 ( TMEMD1 ) ,.TMEMA6 ( TMEMA6 )
 ,.TMEMD0 ( TMEMD0 ) ,.TMEMA5 ( TMEMA5 ) ,.TMEMA4 ( TMEMA4 ) ,.TMEMA3 ( TMEMA3 ) ,.TMEMA2 ( TMEMA2 ) ,.TMEMA1 ( TMEMA1 )
 ,.TMEMA0 ( TMEMA0 ) ,.TMEMCS_B ( TMEMCS_B ) ,.TMEMRD_B ( TMEMRD_B ) ,.TMEMWR_B ( TMEMWR_B ) ,.TMEMCLK2 ( TMEMCLK2 ) ,.TMEMCLK1 ( TMEMCLK1 )
 ,.TMEMCLK0 ( TMEMCLK0 ) ,.TMEMD107 ( TMEMD107 ) ,.TMEMD106 ( TMEMD106 ) ,.TMEMD105 ( TMEMD105 ) ,.TMEMD104 ( TMEMD104 ) ,.TMEMD103 ( TMEMD103 )
 ,.TMEMD102 ( TMEMD102 ) ,.TMEMD101 ( TMEMD101 ) ,.TMEMD100 ( TMEMD100 ) ,.TMEMD99 ( TMEMD99 ) ,.TMEMD98 ( TMEMD98 ) ,.TMEMD97 ( TMEMD97 )
 ,.TMEMD89 ( TMEMD89 ) ,.TMEMD96 ( TMEMD96 ) ,.TMEMD88 ( TMEMD88 ) ,.TMEMD95 ( TMEMD95 ) ,.TMEMD87 ( TMEMD87 ) ,.TMEMD79 ( TMEMD79 )
 ,.TMEMD94 ( TMEMD94 ) ,.TMEMD86 ( TMEMD86 ) ,.TMEMD78 ( TMEMD78 ) ,.TMEMD93 ( TMEMD93 ) ,.TMEMD85 ( TMEMD85 ) ,.TMEMD77 ( TMEMD77 )
 ,.TMEMD69 ( TMEMD69 ) ,.TMEMD92 ( TMEMD92 ) ,.TMEMD84 ( TMEMD84 ) ,.TMEMD76 ( TMEMD76 ) ,.TMEMD68 ( TMEMD68 ) ,.TMEMD91 ( TMEMD91 )
 ,.TMEMD83 ( TMEMD83 ) ,.TMEMD75 ( TMEMD75 ) ,.TMEMD67 ( TMEMD67 ) ,.TMEMD59 ( TMEMD59 ) ,.TMEMD90 ( TMEMD90 ) ,.TMEMD82 ( TMEMD82 )
 ,.TMEMD74 ( TMEMD74 ) ,.TMEMD66 ( TMEMD66 ) ,.TMEMD58 ( TMEMD58 ) ,.TMEMD81 ( TMEMD81 ) ,.TMEMD73 ( TMEMD73 ) ,.TMEMD65 ( TMEMD65 )
 ,.TMEMD57 ( TMEMD57 ) ,.TMEMD49 ( TMEMD49 ) ,.TMEMD80 ( TMEMD80 ) ,.TMEMD72 ( TMEMD72 ) ,.TMEMD64 ( TMEMD64 ) ,.TMEMD56 ( TMEMD56 )
 ,.TMEMD48 ( TMEMD48 ) ,.TMEMD71 ( TMEMD71 ) ,.TMEMD63 ( TMEMD63 ) ,.TMEMD55 ( TMEMD55 ) ,.TMEMD47 ( TMEMD47 ) ,.TMEMD39 ( TMEMD39 )
 ,.TMEMD70 ( TMEMD70 ) ,.TMEMD62 ( TMEMD62 ) ,.TMEMD54 ( TMEMD54 ) ,.TMEMD46 ( TMEMD46 ) ,.TMEMD38 ( TMEMD38 ) ,.TMEMD61 ( TMEMD61 )
 ,.TMEMD53 ( TMEMD53 ) ,.TMEMD45 ( TMEMD45 ) ,.TMEMD37 ( TMEMD37 ) ,.TMEMD29 ( TMEMD29 ) ,.TMEMD60 ( TMEMD60 ) ,.TMEMD52 ( TMEMD52 )
 ,.TMEMD44 ( TMEMD44 ) ,.TMEMD36 ( TMEMD36 ) ,.TMEMD28 ( TMEMD28 ) ,.TMEMD51 ( TMEMD51 ) ,.TMEMD43 ( TMEMD43 ) ,.TMEMD35 ( TMEMD35 )
 ,.TMEMD27 ( TMEMD27 ) ,.TMEMD19 ( TMEMD19 ) ,.TMEMD50 ( TMEMD50 ) ,.TMEMD42 ( TMEMD42 ) ,.TMEMD34 ( TMEMD34 ) ,.TMEMD26 ( TMEMD26 )
 ,.TMEMD18 ( TMEMD18 ) ,.TMEMD41 ( TMEMD41 ) ,.TMEMD33 ( TMEMD33 ) ,.TMEMD25 ( TMEMD25 ) ,.TMEMD17 ( TMEMD17 ) ,.TMEMD40 ( TMEMD40 )
 ,.TMEMD32 ( TMEMD32 ) ,.TMEMD24 ( TMEMD24 ) ,.TMEMD16 ( TMEMD16 ) ,.TMEMD31 ( TMEMD31 ) ,.TMEMD23 ( TMEMD23 ) ,.TMEMD15 ( TMEMD15 )
 ,.TMEMD30 ( TMEMD30 ) ,.TMEMD22 ( TMEMD22 ) ,.TMEMD14 ( TMEMD14 ) ,.TMEMD21 ( TMEMD21 ) ,.TMEMD13 ( TMEMD13 ) ,.TMEMD20 ( TMEMD20 )
 ,.TMEMD12 ( TMEMD12 ) ,.TMEMD11 ( TMEMD11 ) ,.TMEMD10 ( TMEMD10 ) ,.TMEMD9 ( TMEMD9 ) ,.TMEMD8 ( TMEMD8 ) ,.TMEMD7 ( TMEMD7 )
 ,.TMEMD6 ( TMEMD6 ) ,.TMEMD5 ( TMEMD5 ) ,.TMEMD4 ( TMEMD4 )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/eventv1.v
  EVENTV1 eventv1 (
   .CPURESETB ( CPURSOUTB ) ,.EVD21 ( BRKSNAP2 ) ,.EVD13 ( EVD13 ) ,.EVD05 ( EVD05 ) ,.EVD20 ( BRKSNAP1 ) ,.EVD12 ( EVD12 ) ,.EVD04 ( EVD04 )
 ,.EVD19 ( BRKSNAP0 ) ,.EVD18 ( BRKEDMM3 ) ,.EVD17 ( BRKEDMM2 ) ,.EVD09 ( EVD09 ) ,.EVD16 ( BRKEDMM1 ) ,.EVD08 ( EVD08 )
 ,.EVD15 ( BRKEDMM0 ) ,.EVD07 ( EVD07 ) ,.ICEDO31 ( ICEDOK31 ) ,.ICEDO23 ( ICEDOK23 ) ,.ICEDO15 ( ICEDOK15 ) ,.ICEDO30 ( ICEDOK30 )
 ,.ICEDO22 ( ICEDOK22 ) ,.ICEDO14 ( ICEDOK14 ) ,.ICEDO29 ( ICEDOK29 ) ,.ICEDO28 ( ICEDOK28 ) ,.ICEDO27 ( ICEDOK27 ) ,.ICEDO19 ( ICEDOK19 )
 ,.ICEDO26 ( ICEDOK26 ) ,.ICEDO18 ( ICEDOK18 ) ,.ICEDO25 ( ICEDOK25 ) ,.ICEDO17 ( ICEDOK17 ) ,.ICEDO24 ( ICEDOK24 ) ,.ICEDO16 ( ICEDOK16 )
 ,.ICEDO21 ( ICEDOK21 ) ,.ICEDO13 ( ICEDOK13 ) ,.ICEDO20 ( ICEDOK20 ) ,.ICEDO12 ( ICEDOK12 ) ,.ICEDO11 ( ICEDOK11 ) ,.ICEDO10 ( ICEDOK10 )
 ,.ICEDO9 ( ICEDOK9 ) ,.ICEDO8 ( ICEDOK8 ) ,.ICEDO7 ( ICEDOK7 ) ,.ICEDO6 ( ICEDOK6 ) ,.ICEDO5 ( ICEDOK5 ) ,.ICEDO4 ( ICEDOK4 )
 ,.ICEDO3 ( ICEDOK3 ) ,.ICEDO2 ( ICEDOK2 ) ,.ICEDO1 ( ICEDOK1 ) ,.ICEDO0 ( ICEDOK0 ) ,.ICEIFA31 ( ICEIFA31 ) ,.ICEIFA23 ( ICEIFA23 )
 ,.ICEIFA15 ( ICEIFA15 ) ,.ICEIFA30 ( ICEIFA30 ) ,.ICEIFA22 ( ICEIFA22 ) ,.ICEIFA14 ( ICEIFA14 ) ,.ICEIFA29 ( ICEIFA29 ) ,.ICEIFA28 ( ICEIFA28 )
 ,.ICEIFA27 ( ICEIFA27 ) ,.ICEIFA19 ( ICEIFA19 ) ,.ICEIFA26 ( ICEIFA26 ) ,.ICEIFA18 ( ICEIFA18 ) ,.ICEIFA25 ( ICEIFA25 ) ,.ICEIFA17 ( ICEIFA17 )
 ,.ICEIFA24 ( ICEIFA24 ) ,.ICEIFA16 ( ICEIFA16 ) ,.ICEIFA21 ( ICEIFA21 ) ,.ICEIFA13 ( ICEIFA13 ) ,.ICEIFA20 ( ICEIFA20 ) ,.ICEIFA12 ( ICEIFA12 )
 ,.ICEIFA11 ( ICEIFA11 ) ,.ICEIFA10 ( ICEIFA10 ) ,.ICEIFA9 ( ICEIFA9 ) ,.ICEIFA8 ( ICEIFA8 ) ,.ICEIFA7 ( ICEIFA7 ) ,.ICEIFA6 ( ICEIFA6 )
 ,.ICEIFA5 ( ICEIFA5 ) ,.ICEIFA4 ( ICEIFA4 ) ,.ICEIFA3 ( ICEIFA3 ) ,.ICEIFA2 ( ICEIFA2 ) ,.ICEDI19 ( ICEDI19 ) ,.ICEDI18 ( ICEDI18 )
 ,.ICEDI17 ( ICEDI17 ) ,.ICEDI16 ( ICEDI16 ) ,.ICEDI15 ( ICEDI15 ) ,.ICEDI14 ( ICEDI14 ) ,.ICEDI13 ( ICEDI13 ) ,.ICEDI12 ( ICEDI12 )
 ,.ICEDI11 ( ICEDI11 ) ,.ICEDI10 ( ICEDI10 ) ,.ICEDI9 ( ICEDI9 ) ,.ICEDI8 ( ICEDI8 ) ,.ICEDI7 ( ICEDI7 ) ,.ICEDI6 ( ICEDI6 )
 ,.ICEDI5 ( ICEDI5 ) ,.ICEDI4 ( ICEDI4 ) ,.ICEDI3 ( ICEDI3 ) ,.ICEDI2 ( ICEDI2 ) ,.ICEDI1 ( ICEDI1 ) ,.ICEDI0 ( ICEDI0 )
 ,.ICEWR ( ICEWR ) ,.PC19 ( PC19 ) ,.PC18 ( PC18 ) ,.PC17 ( PC17 ) ,.PC16 ( PC16 ) ,.PC15 ( PC15 )
 ,.PC14 ( PC14 ) ,.PC13 ( PC13 ) ,.PC12 ( PC12 ) ,.PC11 ( PC11 ) ,.PC10 ( PC10 ) ,.PC9 ( PC9 )
 ,.PC8 ( PC8 ) ,.PC7 ( PC7 ) ,.PC6 ( PC6 ) ,.PC5 ( PC5 ) ,.PC4 ( PC4 ) ,.PC3 ( PC3 )
 ,.PC2 ( PC2 ) ,.PC1 ( PC1 ) ,.PC0 ( PC0 ) ,.MA15 ( MA15 ) ,.MA14 ( MA14 ) ,.MA13 ( MA13 )
 ,.MA12 ( MA12 ) ,.MA11 ( MA11 ) ,.MA10 ( MA10 ) ,.MA9 ( MA9 ) ,.MA8 ( MA8 ) ,.MA7 ( MA7 )
 ,.MA6 ( MA6 ) ,.MA5 ( MA5 ) ,.MA4 ( MA4 ) ,.MA3 ( MA3 ) ,.MA2 ( MA2 ) ,.MA1 ( MA1 )
 ,.MA0 ( MA0 ) ,.IMDR15 ( IMDR15 ) ,.IMDR14 ( IMDR14 ) ,.IMDR13 ( IMDR13 ) ,.IMDR12 ( IMDR12 ) ,.IMDR11 ( IMDR11 )
 ,.IMDR10 ( IMDR10 ) ,.FLREAD ( FLREAD ) ,.IMDR9 ( IMDR9 ) ,.IMDR8 ( IMDR8 ) ,.IMDR7 ( IMDR7 ) ,.MDW15 ( MDW15 )
 ,.IMDR6 ( IMDR6 ) ,.MDW14 ( MDW14 ) ,.IMDR5 ( IMDR5 ) ,.MDW13 ( MDW13 ) ,.IMDR4 ( IMDR4 ) ,.MDW12 ( MDW12 )
 ,.IMDR3 ( IMDR3 ) ,.MDW11 ( MDW11 ) ,.IMDR2 ( IMDR2 ) ,.MDW10 ( MDW10 ) ,.IMDR1 ( IMDR1 ) ,.IMDR0 ( IMDR0 )
 ,.MDW9 ( MDW9 ) ,.MDW8 ( MDW8 ) ,.MDW7 ( MDW7 ) ,.MDW6 ( MDW6 ) ,.MDW5 ( MDW5 ) ,.MDW4 ( MDW4 )
 ,.MDW3 ( MDW3 ) ,.MDW2 ( MDW2 ) ,.MDW1 ( MDW1 ) ,.MDW0 ( MDW0 ) ,.CPURD ( CPURD ) ,.CPUWR ( CPUWR )
 ,.WDOP ( WDOP ) ,.BASECK ( BASECK ) ,.SYSRSOUTB ( SYSRSOUTB ) ,.TRCON ( TRCON ) ,.TRCMD ( TRCMD ) ,.SELFMODEDBG ( SELFMODEDBG )
 ,.SVMOD ( SVMOD ) ,.SVMODUSER ( SVMODUSER ) ,.STAGEADR1 ( STAGEADR1 ) ,.STAGEADR0 ( STAGEADR0 ) ,.FLREADB3 ( FLREADB3 ) ,.FLREADB2 ( FLREADB2 )
 ,.FLREADB1 ( FLREADB1 ) ,.FLREADB0 ( FLREADB0 ) ,.EROMPD31 ( EROMPD31 ) ,.EROMPD23 ( EROMPD23 ) ,.EROMPD15 ( EROMPD15 ) ,.EROMPD30 ( EROMPD30 )
 ,.EROMPD22 ( EROMPD22 ) ,.EROMPD14 ( EROMPD14 ) ,.EROMPD29 ( EROMPD29 ) ,.EROMPD28 ( EROMPD28 ) ,.EROMPD27 ( EROMPD27 ) ,.EROMPD19 ( EROMPD19 )
 ,.EROMPD26 ( EROMPD26 ) ,.EROMPD18 ( EROMPD18 ) ,.EROMPD25 ( EROMPD25 ) ,.EROMPD17 ( EROMPD17 ) ,.EROMPD24 ( EROMPD24 ) ,.EROMPD16 ( EROMPD16 )
 ,.EROMPD21 ( EROMPD21 ) ,.EROMPD13 ( EROMPD13 ) ,.EROMPD20 ( EROMPD20 ) ,.EROMPD12 ( EROMPD12 ) ,.EROMPD11 ( EROMPD11 ) ,.EROMPD10 ( EROMPD10 )
 ,.EROMPD9 ( EROMPD9 ) ,.EROMPD8 ( EROMPD8 ) ,.EROMPD7 ( EROMPD7 ) ,.EROMPD6 ( EROMPD6 ) ,.EROMPD5 ( EROMPD5 ) ,.EROMPD4 ( EROMPD4 )
 ,.EROMPD3 ( EROMPD3 ) ,.EROMPD2 ( EROMPD2 ) ,.EROMPD1 ( EROMPD1 ) ,.EROMPD0 ( EROMPD0 ) ,.PCWAITF ( PCWAITF ) ,.WAITEXM ( WAITEXM )
 ,.OCDWAIT ( OCDWAIT ) ,.SKIPEXE ( SKIPEXE ) ,.FCHRAM ( FCHRAM ) ,.CPUMASK ( CPUMASK ) ,.INTACK ( INTACK ) ,.DMAACK ( DMAACK )
 ,.EXMA3 ( EXMA3 ) ,.EXMA2 ( EXMA2 ) ,.EXMA1 ( EXMA1 ) ,.EXMA0 ( EXMA0 ) ,.SELEXMPC ( SELEXMPC ) ,.SELRAMPC ( SELRAMPC )
 ,.SELROMPC ( SELROMPC ) ,.SELBRAMPC ( SELBRAMPC ) ,.SELBFAPC ( SELBFAPC ) ,.BRKEVTL1 ( BRKEVTL1 ) ,.BRKEVTL0 ( BRKEVTL0 ) ,.BRKEVTA7 ( BRKEVTA7 )
 ,.BRKEVTA6 ( BRKEVTA6 ) ,.BRKEVTA5 ( BRKEVTA5 ) ,.BRKEVTA4 ( BRKEVTA4 ) ,.BRKEVTA3 ( BRKEVTA3 ) ,.BRKEVTA2 ( BRKEVTA2 ) ,.BRKEVTA1 ( BRKEVTA1 )
 ,.BRKEVTA0 ( BRKEVTA0 ) ,.BRKEVTF7 ( BRKEVTF7 ) ,.BRKEVTF6 ( BRKEVTF6 ) ,.BRKEVTF5 ( BRKEVTF5 ) ,.BRKEVTF4 ( BRKEVTF4 ) ,.BRKEVTF3 ( BRKEVTF3 )
 ,.BRKEVTF2 ( BRKEVTF2 ) ,.BRKEVTF1 ( BRKEVTF1 ) ,.BRKEVTF0 ( BRKEVTF0 ) ,.EVD14 ( EVD14 ) ,.EVD06 ( EVD06 ) ,.EVD11 ( EVD11 )
 ,.EVD03 ( EVD03 ) ,.EVD10 ( EVD10 ) ,.EVD02 ( EVD02 ) ,.EVD01 ( EVD01 )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/failsafev1.v
  FAILSAFEV1 failsafe (
   .CK60MHZ ( CLK30MHZ_GB ) ,.CPURESETB ( CPURSOUTB ) ,.ICEDO31 ( ICEDOH31 ) ,.ICEDO23 ( ICEDOH23 ) ,.ICEDO15 ( ICEDOH15 ) ,.ICEDO30 ( ICEDOH30 ) ,.ICEDO22 ( ICEDOH22 )
 ,.ICEDO14 ( ICEDOH14 ) ,.ICEDO29 ( ICEDOH29 ) ,.ICEDO28 ( ICEDOH28 ) ,.ICEDO27 ( ICEDOH27 ) ,.ICEDO19 ( ICEDOH19 ) ,.ICEDO26 ( ICEDOH26 )
 ,.ICEDO18 ( ICEDOH18 ) ,.ICEDO25 ( ICEDOH25 ) ,.ICEDO17 ( ICEDOH17 ) ,.ICEDO24 ( ICEDOH24 ) ,.ICEDO16 ( ICEDOH16 ) ,.ICEDO21 ( ICEDOH21 )
 ,.ICEDO13 ( ICEDOH13 ) ,.ICEDO20 ( ICEDOH20 ) ,.ICEDO12 ( ICEDOH12 ) ,.ICEDO11 ( ICEDOH11 ) ,.ICEDO10 ( ICEDOH10 ) ,.ICEDO9 ( ICEDOH9 )
 ,.ICEDO8 ( ICEDOH8 ) ,.ICEDO7 ( ICEDOH7 ) ,.ICEDO6 ( ICEDOH6 ) ,.ICEDO5 ( ICEDOH5 ) ,.ICEDO4 ( ICEDOH4 ) ,.ICEDO3 ( ICEDOH3 )
 ,.ICEDO2 ( ICEDOH2 ) ,.ICEDO1 ( ICEDOH1 ) ,.ICEDO0 ( ICEDOH0 ) ,.ICEIFA31 ( ICEIFA31 ) ,.ICEIFA23 ( ICEIFA23 ) ,.ICEIFA15 ( ICEIFA15 )
 ,.ICEIFA30 ( ICEIFA30 ) ,.ICEIFA22 ( ICEIFA22 ) ,.ICEIFA14 ( ICEIFA14 ) ,.ICEIFA29 ( ICEIFA29 ) ,.ICEIFA28 ( ICEIFA28 ) ,.ICEIFA27 ( ICEIFA27 )
 ,.ICEIFA19 ( ICEIFA19 ) ,.ICEIFA26 ( ICEIFA26 ) ,.ICEIFA18 ( ICEIFA18 ) ,.ICEIFA25 ( ICEIFA25 ) ,.ICEIFA17 ( ICEIFA17 ) ,.ICEIFA24 ( ICEIFA24 )
 ,.ICEIFA16 ( ICEIFA16 ) ,.ICEIFA21 ( ICEIFA21 ) ,.ICEIFA13 ( ICEIFA13 ) ,.ICEIFA20 ( ICEIFA20 ) ,.ICEIFA12 ( ICEIFA12 ) ,.ICEIFA11 ( ICEIFA11 )
 ,.ICEIFA10 ( ICEIFA10 ) ,.ICEIFA9 ( ICEIFA9 ) ,.ICEIFA8 ( ICEIFA8 ) ,.ICEIFA7 ( ICEIFA7 ) ,.ICEIFA6 ( ICEIFA6 ) ,.ICEIFA5 ( ICEIFA5 )
 ,.ICEIFA4 ( ICEIFA4 ) ,.ICEIFA3 ( ICEIFA3 ) ,.ICEIFA2 ( ICEIFA2 ) ,.ICEDI31 ( ICEDI31 ) ,.ICEDI23 ( ICEDI23 ) ,.ICEDI15 ( ICEDI15 )
 ,.ICEDI30 ( ICEDI30 ) ,.ICEDI22 ( ICEDI22 ) ,.ICEDI14 ( ICEDI14 ) ,.ICEDI29 ( ICEDI29 ) ,.ICEDI28 ( ICEDI28 ) ,.ICEDI27 ( ICEDI27 )
 ,.ICEDI19 ( ICEDI19 ) ,.ICEDI26 ( ICEDI26 ) ,.ICEDI18 ( ICEDI18 ) ,.ICEDI25 ( ICEDI25 ) ,.ICEDI17 ( ICEDI17 ) ,.ICEDI24 ( ICEDI24 )
 ,.ICEDI16 ( ICEDI16 ) ,.ICEDI21 ( ICEDI21 ) ,.ICEDI13 ( ICEDI13 ) ,.ICEDI20 ( ICEDI20 ) ,.ICEDI12 ( ICEDI12 ) ,.ICEDI11 ( ICEDI11 )
 ,.ICEDI10 ( ICEDI10 ) ,.ICEDI9 ( ICEDI9 ) ,.ICEDI8 ( ICEDI8 ) ,.ICEDI7 ( ICEDI7 ) ,.ICEDI6 ( ICEDI6 ) ,.ICEDI5 ( ICEDI5 )
 ,.ICEDI4 ( ICEDI4 ) ,.ICEDI3 ( ICEDI3 ) ,.ICEDI2 ( ICEDI2 ) ,.ICEDI1 ( ICEDI1 ) ,.ICEDI0 ( ICEDI0 ) ,.ICEWR ( ICEWR )
 ,.PC19 ( PC19 ) ,.PC18 ( PC18 ) ,.PC17 ( PC17 ) ,.PC16 ( PC16 ) ,.PC15 ( PC15 ) ,.PC14 ( PC14 )
 ,.PC13 ( PC13 ) ,.PC12 ( PC12 ) ,.PC11 ( PC11 ) ,.PC10 ( PC10 ) ,.PC9 ( PC9 ) ,.PC8 ( PC8 )
 ,.PC7 ( PC7 ) ,.PC6 ( PC6 ) ,.PC5 ( PC5 ) ,.PC4 ( PC4 ) ,.PC3 ( PC3 ) ,.PC2 ( PC2 )
 ,.PC1 ( PC1 ) ,.PC0 ( PC0 ) ,.FLMA15 ( FLMA15 ) ,.FLMA14 ( FLMA14 ) ,.FLMA13 ( FLMA13 ) ,.FLMA12 ( FLMA12 )
 ,.FLMA11 ( FLMA11 ) ,.FLMA10 ( FLMA10 ) ,.FLMA9 ( FLMA9 ) ,.FLMA8 ( FLMA8 ) ,.FLMA7 ( FLMA7 ) ,.FLMA6 ( FLMA6 )
 ,.FLMA5 ( FLMA5 ) ,.FLMA4 ( FLMA4 ) ,.FLMA3 ( FLMA3 ) ,.FLMA2 ( FLMA2 ) ,.FLMA1 ( FLMA1 ) ,.FLMA0 ( FLMA0 )
 ,.EXMA3 ( EXMA3 ) ,.EXMA2 ( EXMA2 ) ,.EXMA1 ( EXMA1 ) ,.EXMA0 ( EXMA0 ) ,.BASECK ( BASECK ) ,.CPURD ( CPURD )
 ,.CPUWR ( CPUWR ) ,.WDOP ( WDOP ) ,.SVMOD ( SVMOD ) ,.MAAOUT ( MAAOUT ) ,.STAGEADR1 ( STAGEADR1 ) ,.STAGEADR0 ( STAGEADR0 )
 ,.PCWAITF ( PCWAITF ) ,.SKIPEXE ( SKIPEXE ) ,.FCHRAM ( FCHRAM ) ,.ALT1 ( ALT1 ) ,.IDPOP ( IDPOP ) ,.SPINC ( SPINC )
 ,.SPDEC ( SPDEC ) ,.SPREL ( SPREL ) ,.CPUMISAL ( CPUMISAL ) ,.SYSRSOUTB ( SYSRSOUTB ) ,.PERISVIB ( PERISVIB ) ,.SELFMODE ( SELFMODE )
 ,.BRAMEN ( BRAMEN ) ,.BFAEN ( BFAEN ) ,.INTACK ( INTACK ) ,.DMAACK ( DMAACK ) ,.WAITEXM ( WAITEXM ) ,.OCDWAIT ( OCDWAIT )
 ,.SOFTBRK ( SOFTBRK ) ,.FLSIZE3 ( FLSIZE3 ) ,.FLSIZE2 ( FLSIZE2 ) ,.FLSIZE1 ( FLSIZE1 ) ,.FLSIZE0 ( FLSIZE0 ) ,.RAMSIZE7 ( RAMSIZE7 )
 ,.RAMSIZE6 ( RAMSIZE6 ) ,.RAMSIZE5 ( RAMSIZE5 ) ,.RAMSIZE4 ( RAMSIZE4 ) ,.RAMSIZE3 ( RAMSIZE3 ) ,.RAMSIZE2 ( RAMSIZE2 ) ,.RAMSIZE1 ( RAMSIZE1 )
 ,.RAMSIZE0 ( RAMSIZE0 ) ,.BFSIZE3 ( BFSIZE3 ) ,.BFSIZE2 ( BFSIZE2 ) ,.BFSIZE1 ( BFSIZE1 ) ,.BFSIZE0 ( BFSIZE0 ) ,.BMSIZE3 ( BMSIZE3 )
 ,.BMSIZE2 ( BMSIZE2 ) ,.BMSIZE1 ( BMSIZE1 ) ,.BMSIZE0 ( BMSIZE0 ) ,.DFSIZE1 ( DFSIZE1 ) ,.DFSIZE0 ( DFSIZE0 ) ,.BRKFAIL0 ( BRKFAIL0 )
 ,.BRKFAIL1 ( BRKFAIL1 ) ,.BRKFAIL2 ( BRKFAIL2 ) ,.BRKFAIL3 ( BRKFAIL3 ) ,.BRKFAIL4 ( BRKFAIL4 ) ,.BRKFAIL5 ( BRKFAIL5 ) ,.BRKFAIL6 ( BRKFAIL6 )
 ,.BRKFAIL7 ( BRKFAIL7 ) ,.BRKFAIL8 ( BRKFAIL8 ) ,.BRKFAIL9 ( BRKFAIL9 ) ,.BRKFAIL10 ( BRKFAIL10 ) ,.BRKFAIL11 ( BRKFAIL11 ) ,.BRKFAIL13 ( BRKFAIL13 )
 ,.BRKFAIL15 ( BRKFAIL15 ) ,.FAILMK12 ( FAILMK12 ) ,.EXMAPOUT ( EXMAPOUT ) ,.SELEXMPC ( SELEXMPC ) ,.SELRAMPC ( SELRAMPC ) ,.SELROMPC ( SELROMPC )
 ,.SELBRAMPC ( SELBRAMPC ) ,.SELBFAPC ( SELBFAPC ) ,.SELRAMMA ( SELRAMMA ) ,.SELDFADMA ( SELDFADMA )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/pseudoemu.v
  PSEUDOEMU pseudoemu (
   .ICEDO31 ( ICEDOQ31 ) ,.ICEDO23 ( ICEDOQ23 ) ,.ICEDO15 ( ICEDOQ15 ) ,.ICEDO30 ( ICEDOQ30 ) ,.ICEDO22 ( ICEDOQ22 ) ,.ICEDO14 ( ICEDOQ14 ) ,.ICEDO29 ( ICEDOQ29 )
 ,.ICEDO28 ( ICEDOQ28 ) ,.ICEDO27 ( ICEDOQ27 ) ,.ICEDO19 ( ICEDOQ19 ) ,.ICEDO26 ( ICEDOQ26 ) ,.ICEDO18 ( ICEDOQ18 ) ,.ICEDO25 ( ICEDOQ25 )
 ,.ICEDO17 ( ICEDOQ17 ) ,.ICEDO24 ( ICEDOQ24 ) ,.ICEDO16 ( ICEDOQ16 ) ,.ICEDO21 ( ICEDOQ21 ) ,.ICEDO13 ( ICEDOQ13 ) ,.ICEDO20 ( ICEDOQ20 )
 ,.ICEDO12 ( ICEDOQ12 ) ,.ICEDO11 ( ICEDOQ11 ) ,.ICEDO10 ( ICEDOQ10 ) ,.ICEDO9 ( ICEDOQ9 ) ,.ICEDO8 ( ICEDOQ8 ) ,.ICEDO7 ( ICEDOQ7 )
 ,.ICEDO6 ( ICEDOQ6 ) ,.ICEDO5 ( ICEDOQ5 ) ,.ICEDO4 ( ICEDOQ4 ) ,.ICEDO3 ( ICEDOQ3 ) ,.ICEDO2 ( ICEDOQ2 ) ,.ICEDO1 ( ICEDOQ1 )
 ,.ICEDO0 ( ICEDOQ0 ) ,.ICEIFA31 ( ICEIFA31 ) ,.ICEIFA23 ( ICEIFA23 ) ,.ICEIFA15 ( ICEIFA15 ) ,.ICEIFA30 ( ICEIFA30 ) ,.ICEIFA22 ( ICEIFA22 )
 ,.ICEIFA14 ( ICEIFA14 ) ,.ICEIFA29 ( ICEIFA29 ) ,.ICEIFA28 ( ICEIFA28 ) ,.ICEIFA27 ( ICEIFA27 ) ,.ICEIFA19 ( ICEIFA19 ) ,.ICEIFA26 ( ICEIFA26 )
 ,.ICEIFA18 ( ICEIFA18 ) ,.ICEIFA25 ( ICEIFA25 ) ,.ICEIFA17 ( ICEIFA17 ) ,.ICEIFA24 ( ICEIFA24 ) ,.ICEIFA16 ( ICEIFA16 ) ,.ICEIFA21 ( ICEIFA21 )
 ,.ICEIFA13 ( ICEIFA13 ) ,.ICEIFA20 ( ICEIFA20 ) ,.ICEIFA12 ( ICEIFA12 ) ,.ICEIFA11 ( ICEIFA11 ) ,.ICEIFA10 ( ICEIFA10 ) ,.ICEIFA9 ( ICEIFA9 )
 ,.ICEIFA8 ( ICEIFA8 ) ,.ICEIFA7 ( ICEIFA7 ) ,.ICEIFA6 ( ICEIFA6 ) ,.ICEIFA5 ( ICEIFA5 ) ,.ICEIFA4 ( ICEIFA4 ) ,.ICEIFA3 ( ICEIFA3 )
 ,.ICEIFA2 ( ICEIFA2 ) ,.ICEIFA1 ( ICEIFA1 ) ,.ICEIFA0 ( ICEIFA0 ) ,.ICEDI15 ( ICEDI15 ) ,.ICEDI14 ( ICEDI14 ) ,.ICEDI13 ( ICEDI13 )
 ,.ICEDI12 ( ICEDI12 ) ,.ICEDI11 ( ICEDI11 ) ,.ICEDI10 ( ICEDI10 ) ,.ICEDI9 ( ICEDI9 ) ,.ICEDI8 ( ICEDI8 ) ,.ICEDI7 ( ICEDI7 )
 ,.ICEDI6 ( ICEDI6 ) ,.ICEDI5 ( ICEDI5 ) ,.ICEDI4 ( ICEDI4 ) ,.ICEDI3 ( ICEDI3 ) ,.ICEDI2 ( ICEDI2 ) ,.ICEDI1 ( ICEDI1 )
 ,.ICEDI0 ( ICEDI0 ) ,.ICEWR ( ICEWR ) ,.PSEUDOON31 ( PSEUDOON31 ) ,.PSEUDOON23 ( PSEUDOON23 ) ,.PSEUDOON15 ( PSEUDOON15 ) ,.PSEUDOON30 ( PSEUDOON30 )
 ,.PSEUDOON22 ( PSEUDOON22 ) ,.PSEUDOON14 ( PSEUDOON14 ) ,.PSEUDOON29 ( PSEUDOON29 ) ,.PSEUDOON28 ( PSEUDOON28 ) ,.PSEUDOON27 ( PSEUDOON27 ) ,.PSEUDOON19 ( PSEUDOON19 )
 ,.PSEUDOON26 ( PSEUDOON26 ) ,.PSEUDOON18 ( PSEUDOON18 ) ,.PSEUDOON25 ( PSEUDOON25 ) ,.PSEUDOON17 ( PSEUDOON17 ) ,.PSEUDOON24 ( PSEUDOON24 ) ,.PSEUDOON16 ( PSEUDOON16 )
 ,.PSEUDOON21 ( PSEUDOON21 ) ,.PSEUDOON13 ( PSEUDOON13 ) ,.PSEUDOON20 ( PSEUDOON20 ) ,.PSEUDOON12 ( PSEUDOON12 ) ,.PSEUDOON11 ( PSEUDOON11 ) ,.PSEUDOON10 ( PSEUDOON10 )
 ,.PSEUDOON9 ( PSEUDOON9 ) ,.PSEUDOON8 ( PSEUDOON8 ) ,.PSEUDOON7 ( PSEUDOON7 ) ,.PSEUDOON6 ( PSEUDOON6 ) ,.PSEUDOON5 ( PSEUDOON5 ) ,.PSEUDOON4 ( PSEUDOON4 )
 ,.PSEUDOON3 ( PSEUDOON3 ) ,.PSEUDOON2 ( PSEUDOON2 ) ,.PSEUDOON1 ( PSEUDOON1 ) ,.PSEUDOON0 ( PSEUDOON0 ) ,.PSEUDORES ( PSEUDORES ) ,.SYSRSOUTB ( SYSRSOUTB )
 ,.SVMOD ( SVMOD ) ,.PSEUDOANI09 ( PSEUDOANI09 ) ,.PSEUDOANI17 ( PSEUDOANI17 ) ,.PSEUDOANI08 ( PSEUDOANI08 ) ,.PSEUDOANI16 ( PSEUDOANI16 ) ,.PSEUDOANI07 ( PSEUDOANI07 )
 ,.PSEUDOANI15 ( PSEUDOANI15 ) ,.PSEUDOANI06 ( PSEUDOANI06 ) ,.PSEUDOANI14 ( PSEUDOANI14 ) ,.PSEUDOANI05 ( PSEUDOANI05 ) ,.PSEUDOANI13 ( PSEUDOANI13 ) ,.PSEUDOANI04 ( PSEUDOANI04 )
 ,.PSEUDOANI12 ( PSEUDOANI12 ) ,.PSEUDOANI03 ( PSEUDOANI03 ) ,.PSEUDOANI11 ( PSEUDOANI11 ) ,.PSEUDOANI02 ( PSEUDOANI02 ) ,.PSEUDOANI10 ( PSEUDOANI10 ) ,.PSEUDOANI01 ( PSEUDOANI01 )
 ,.PSEUDOANI00 ( PSEUDOANI00 ) ,.PSEUDOANI19 ( PSEUDOANI19 ) ,.PSEUDOANI18 ( PSEUDOANI18 )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/status.v
  STATUS status (
   .CPURESETB ( CPURSOUTB ) ,.TRESET_B ( TARRESB ) ,.TCCONNECT_B ( ETCCONNECT_B ) ,.EACONNECT_B ( EEACONNECT_B ) ,.TVDDON ( ETVDDON ) ,.TVDDSEL ( ETVDDSEL ) ,.LEDTVDD_B ( ELEDTVDD_B )
 ,.LEDCLOCK_B ( ELEDCLOCK_B ) ,.LEDRUN_B ( ELEDRUN_B ) ,.LEDRESET_B ( ELEDRESET_B ) ,.LEDSTANDBY_B ( ELEDSTANDBY_B ) ,.LEDWAIT_B ( ELEDWAIT_B ) ,.CK60MHZ ( CLK60MHZ )
 ,.TBTSELOUT ( SWAP ) ,.ICEDO31 ( ICEDOJ31 ) ,.ICEDO23 ( ICEDOJ23 ) ,.ICEDO15 ( ICEDOJ15 ) ,.ICEDO30 ( ICEDOJ30 ) ,.ICEDO22 ( ICEDOJ22 )
 ,.ICEDO14 ( ICEDOJ14 ) ,.ICEDO29 ( ICEDOJ29 ) ,.ICEDO28 ( ICEDOJ28 ) ,.ICEDO27 ( ICEDOJ27 ) ,.ICEDO19 ( ICEDOJ19 ) ,.ICEDO26 ( ICEDOJ26 )
 ,.ICEDO18 ( ICEDOJ18 ) ,.ICEDO25 ( ICEDOJ25 ) ,.ICEDO17 ( ICEDOJ17 ) ,.ICEDO24 ( ICEDOJ24 ) ,.ICEDO16 ( ICEDOJ16 ) ,.ICEDO21 ( ICEDOJ21 )
 ,.ICEDO13 ( ICEDOJ13 ) ,.ICEDO20 ( ICEDOJ20 ) ,.ICEDO12 ( ICEDOJ12 ) ,.ICEDO11 ( ICEDOJ11 ) ,.ICEDO10 ( ICEDOJ10 ) ,.ICEDO9 ( ICEDOJ9 )
 ,.ICEDO8 ( ICEDOJ8 ) ,.ICEDO7 ( ICEDOJ7 ) ,.ICEDO6 ( ICEDOJ6 ) ,.ICEDO5 ( ICEDOJ5 ) ,.ICEDO4 ( ICEDOJ4 ) ,.ICEDO3 ( ICEDOJ3 )
 ,.ICEDO2 ( ICEDOJ2 ) ,.ICEDO1 ( ICEDOJ1 ) ,.ICEDO0 ( ICEDOJ0 ) ,.BASECK ( BASECK ) ,.SVMOD ( SVMOD ) ,.SVMODUSER ( SVMODUSER )
 ,.ALT1 ( ALT1 ) ,.SELFMODE ( SELFMODE ) ,.HLTST ( HLTST ) ,.STPST ( STPST ) ,.WAITEXM ( WAITEXM ) ,.EVAOSCMCLK ( EVAOSCMCLK )
 ,.CPUSCLK ( CPUSCLK ) ,.CPUTMCLK ( CPUTMCLK ) ,.WDOP ( WDOP ) ,.CPURD ( CPURD ) ,.CPUWR ( CPUWR ) ,.MA15 ( MA15 )
 ,.MA14 ( MA14 ) ,.MA13 ( MA13 ) ,.MA12 ( MA12 ) ,.MA11 ( MA11 ) ,.MA10 ( MA10 ) ,.MA9 ( MA9 )
 ,.MA8 ( MA8 ) ,.MA7 ( MA7 ) ,.MA6 ( MA6 ) ,.MA5 ( MA5 ) ,.MA4 ( MA4 ) ,.MA3 ( MA3 )
 ,.MA2 ( MA2 ) ,.MA1 ( MA1 ) ,.MA0 ( MA0 ) ,.MDW15 ( MDW15 ) ,.MDW14 ( MDW14 ) ,.MDW13 ( MDW13 )
 ,.MDW12 ( MDW12 ) ,.MDW11 ( MDW11 ) ,.MDW10 ( MDW10 ) ,.MDW9 ( MDW9 ) ,.MDW8 ( MDW8 ) ,.MDW7 ( MDW7 )
 ,.MDW6 ( MDW6 ) ,.MDW5 ( MDW5 ) ,.MDW4 ( MDW4 ) ,.MDW3 ( MDW3 ) ,.MDW2 ( MDW2 ) ,.MDW1 ( MDW1 )
 ,.MDW0 ( MDW0 ) ,.STATEMDR15 ( STATEMDR15 ) ,.STATEMDR14 ( STATEMDR14 ) ,.STATEMDR13 ( STATEMDR13 ) ,.STATEMDR12 ( STATEMDR12 ) ,.STATEMDR11 ( STATEMDR11 )
 ,.STATEMDR10 ( STATEMDR10 ) ,.STATEMDR9 ( STATEMDR9 ) ,.STATEMDR8 ( STATEMDR8 ) ,.STATEMDR7 ( STATEMDR7 ) ,.STATEMDR6 ( STATEMDR6 ) ,.STATEMDR5 ( STATEMDR5 )
 ,.STATEMDR4 ( STATEMDR4 ) ,.STATEMDR3 ( STATEMDR3 ) ,.STATEMDR2 ( STATEMDR2 ) ,.STATEMDR1 ( STATEMDR1 ) ,.STATEMDR0 ( STATEMDR0 ) ,.ICEIFA31 ( ICEIFA31 )
 ,.ICEIFA23 ( ICEIFA23 ) ,.ICEIFA15 ( ICEIFA15 ) ,.ICEIFA30 ( ICEIFA30 ) ,.ICEIFA22 ( ICEIFA22 ) ,.ICEIFA14 ( ICEIFA14 ) ,.ICEIFA29 ( ICEIFA29 )
 ,.ICEIFA28 ( ICEIFA28 ) ,.ICEIFA27 ( ICEIFA27 ) ,.ICEIFA19 ( ICEIFA19 ) ,.ICEIFA26 ( ICEIFA26 ) ,.ICEIFA18 ( ICEIFA18 ) ,.ICEIFA25 ( ICEIFA25 )
 ,.ICEIFA17 ( ICEIFA17 ) ,.ICEIFA24 ( ICEIFA24 ) ,.ICEIFA16 ( ICEIFA16 ) ,.ICEIFA21 ( ICEIFA21 ) ,.ICEIFA13 ( ICEIFA13 ) ,.ICEIFA20 ( ICEIFA20 )
 ,.ICEIFA12 ( ICEIFA12 ) ,.ICEIFA11 ( ICEIFA11 ) ,.ICEIFA10 ( ICEIFA10 ) ,.ICEIFA9 ( ICEIFA9 ) ,.ICEIFA8 ( ICEIFA8 ) ,.ICEIFA7 ( ICEIFA7 )
 ,.ICEIFA6 ( ICEIFA6 ) ,.ICEIFA5 ( ICEIFA5 ) ,.ICEIFA4 ( ICEIFA4 ) ,.ICEIFA3 ( ICEIFA3 ) ,.ICEIFA2 ( ICEIFA2 ) ,.ICEIFA1 ( ICEIFA1 )
 ,.ICEIFA0 ( ICEIFA0 ) ,.ICEDI31 ( ICEDI31 ) ,.ICEDI23 ( ICEDI23 ) ,.ICEDI15 ( ICEDI15 ) ,.ICEDI30 ( ICEDI30 ) ,.ICEDI22 ( ICEDI22 )
 ,.ICEDI14 ( ICEDI14 ) ,.ICEDI29 ( ICEDI29 ) ,.ICEDI28 ( ICEDI28 ) ,.ICEDI27 ( ICEDI27 ) ,.ICEDI19 ( ICEDI19 ) ,.ICEDI26 ( ICEDI26 )
 ,.ICEDI18 ( ICEDI18 ) ,.ICEDI25 ( ICEDI25 ) ,.ICEDI17 ( ICEDI17 ) ,.ICEDI24 ( ICEDI24 ) ,.ICEDI16 ( ICEDI16 ) ,.ICEDI21 ( ICEDI21 )
 ,.ICEDI13 ( ICEDI13 ) ,.ICEDI20 ( ICEDI20 ) ,.ICEDI12 ( ICEDI12 ) ,.ICEDI11 ( ICEDI11 ) ,.ICEDI10 ( ICEDI10 ) ,.ICEDI9 ( ICEDI9 )
 ,.ICEDI8 ( ICEDI8 ) ,.ICEDI7 ( ICEDI7 ) ,.ICEDI6 ( ICEDI6 ) ,.ICEDI5 ( ICEDI5 ) ,.ICEDI4 ( ICEDI4 ) ,.ICEDI3 ( ICEDI3 )
 ,.ICEDI2 ( ICEDI2 ) ,.ICEDI1 ( ICEDI1 ) ,.ICEDI0 ( ICEDI0 ) ,.ICEWR ( ICEWR ) ,.SYSRSOUTB ( SYSRSOUTB )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/coverage.v
  COVERAGE coverage (
   .PA17 ( PA19 ) ,.PA16 ( PA18 ) ,.PA15 ( PA17 ) ,.PA14 ( PA16 ) ,.PA13 ( PA15 ) ,.PA12 ( PA14 ) ,.PA11 ( PA13 )
 ,.PA10 ( PA12 ) ,.PA9 ( PA11 ) ,.PC5 ( PC5 ) ,.PA8 ( PA10 ) ,.PC4 ( PC4 ) ,.PA7 ( PA9 )
 ,.PC3 ( PC3 ) ,.PA6 ( PA8 ) ,.PC2 ( PC2 ) ,.PA5 ( PA7 ) ,.PC1 ( PC1 ) ,.PA4 ( PA6 )
 ,.PC0 ( PC0 ) ,.PA3 ( PA5 ) ,.PA2 ( PA4 ) ,.PA1 ( PA3 ) ,.PA0 ( PA2 ) ,.CPURESETB ( CPURSOUTB )
 ,.CK60MHZ ( CLK60MHZ ) ,.PC19 ( PC19 ) ,.PC18 ( PC18 ) ,.PC17 ( PC17 ) ,.PC16 ( PC16 ) ,.PC15 ( PC15 )
 ,.PC14 ( PC14 ) ,.PC13 ( PC13 ) ,.PC12 ( PC12 ) ,.PC11 ( PC11 ) ,.PC10 ( PC10 ) ,.PC9 ( PC9 )
 ,.PC8 ( PC8 ) ,.PC7 ( PC7 ) ,.PC6 ( PC6 ) ,.ES3 ( EXMA3 ) ,.MA7 ( MA7 ) ,.ES2 ( EXMA2 )
 ,.MA6 ( MA6 ) ,.ES1 ( EXMA1 ) ,.MA5 ( MA5 ) ,.ES0 ( EXMA0 ) ,.MA4 ( MA4 ) ,.ICEDO31 ( ICEDOM31 )
 ,.ICEDO23 ( ICEDOM23 ) ,.ICEDO15 ( ICEDOM15 ) ,.ICEDO30 ( ICEDOM30 ) ,.ICEDO22 ( ICEDOM22 ) ,.ICEDO14 ( ICEDOM14 ) ,.ICEDO29 ( ICEDOM29 )
 ,.ICEDO28 ( ICEDOM28 ) ,.ICEDO27 ( ICEDOM27 ) ,.ICEDO19 ( ICEDOM19 ) ,.ICEDO26 ( ICEDOM26 ) ,.ICEDO18 ( ICEDOM18 ) ,.ICEDO25 ( ICEDOM25 )
 ,.ICEDO17 ( ICEDOM17 ) ,.ICEDO24 ( ICEDOM24 ) ,.ICEDO16 ( ICEDOM16 ) ,.ICEDO21 ( ICEDOM21 ) ,.ICEDO13 ( ICEDOM13 ) ,.ICEDO20 ( ICEDOM20 )
 ,.ICEDO12 ( ICEDOM12 ) ,.ICEDO11 ( ICEDOM11 ) ,.ICEDO10 ( ICEDOM10 ) ,.ICEDO9 ( ICEDOM9 ) ,.ICEDO8 ( ICEDOM8 ) ,.ICEDO7 ( ICEDOM7 )
 ,.ICEDO6 ( ICEDOM6 ) ,.ICEDO5 ( ICEDOM5 ) ,.ICEDO4 ( ICEDOM4 ) ,.ICEDO3 ( ICEDOM3 ) ,.ICEDO2 ( ICEDOM2 ) ,.ICEDO1 ( ICEDOM1 )
 ,.ICEDO0 ( ICEDOM0 ) ,.MA15 ( MA15 ) ,.MA14 ( MA14 ) ,.MA13 ( MA13 ) ,.MA12 ( MA12 ) ,.MA11 ( MA11 )
 ,.MA10 ( MA10 ) ,.MA9 ( MA9 ) ,.MA8 ( MA8 ) ,.MA3 ( MA3 ) ,.MA2 ( MA2 ) ,.MA1 ( MA1 )
 ,.MA0 ( MA0 ) ,.FLREAD ( FLREAD ) ,.FLREADB3 ( FLREADB3 ) ,.FLREADB2 ( FLREADB2 ) ,.FLREADB1 ( FLREADB1 ) ,.FLREADB0 ( FLREADB0 )
 ,.SVMOD ( SVMOD ) ,.SELFMODEDBG ( SELFMODEDBG ) ,.SKIPEXE ( SKIPEXE ) ,.CPUMASK ( CPUMASK ) ,.PCWAITF ( PCWAITF ) ,.STAGEADR0 ( STAGEADR0 )
 ,.STAGEADR1 ( STAGEADR1 ) ,.WAITEXM ( WAITEXM ) ,.SLEXM ( SLEXM ) ,.FCHRAM ( FCHRAM ) ,.WDOP ( WDOP ) ,.CPUWR ( CPUWR )
 ,.CPURD ( CPURD ) ,.INTACK ( INTACK ) ,.DMAACK ( DMAACK ) ,.BASECK ( BASECK ) ,.ICEIFA31 ( ICEIFA31 ) ,.ICEIFA23 ( ICEIFA23 )
 ,.ICEIFA15 ( ICEIFA15 ) ,.ICEIFA30 ( ICEIFA30 ) ,.ICEIFA22 ( ICEIFA22 ) ,.ICEIFA14 ( ICEIFA14 ) ,.ICEIFA29 ( ICEIFA29 ) ,.ICEIFA28 ( ICEIFA28 )
 ,.ICEIFA27 ( ICEIFA27 ) ,.ICEIFA19 ( ICEIFA19 ) ,.ICEIFA26 ( ICEIFA26 ) ,.ICEIFA18 ( ICEIFA18 ) ,.ICEIFA25 ( ICEIFA25 ) ,.ICEIFA17 ( ICEIFA17 )
 ,.ICEIFA24 ( ICEIFA24 ) ,.ICEIFA16 ( ICEIFA16 ) ,.ICEIFA21 ( ICEIFA21 ) ,.ICEIFA13 ( ICEIFA13 ) ,.ICEIFA20 ( ICEIFA20 ) ,.ICEIFA12 ( ICEIFA12 )
 ,.ICEIFA11 ( ICEIFA11 ) ,.ICEIFA10 ( ICEIFA10 ) ,.ICEIFA9 ( ICEIFA9 ) ,.ICEIFA8 ( ICEIFA8 ) ,.ICEIFA7 ( ICEIFA7 ) ,.ICEIFA6 ( ICEIFA6 )
 ,.ICEIFA5 ( ICEIFA5 ) ,.ICEIFA4 ( ICEIFA4 ) ,.ICEIFA3 ( ICEIFA3 ) ,.ICEIFA2 ( ICEIFA2 ) ,.ICEIFA1 ( ICEIFA1 ) ,.ICEIFA0 ( ICEIFA0 )
 ,.ICEDI31 ( ICEDI31 ) ,.ICEDI23 ( ICEDI23 ) ,.ICEDI15 ( ICEDI15 ) ,.ICEDI30 ( ICEDI30 ) ,.ICEDI22 ( ICEDI22 ) ,.ICEDI14 ( ICEDI14 )
 ,.ICEDI29 ( ICEDI29 ) ,.ICEDI28 ( ICEDI28 ) ,.ICEDI27 ( ICEDI27 ) ,.ICEDI19 ( ICEDI19 ) ,.ICEDI26 ( ICEDI26 ) ,.ICEDI18 ( ICEDI18 )
 ,.ICEDI25 ( ICEDI25 ) ,.ICEDI17 ( ICEDI17 ) ,.ICEDI24 ( ICEDI24 ) ,.ICEDI16 ( ICEDI16 ) ,.ICEDI21 ( ICEDI21 ) ,.ICEDI13 ( ICEDI13 )
 ,.ICEDI20 ( ICEDI20 ) ,.ICEDI12 ( ICEDI12 ) ,.ICEDI11 ( ICEDI11 ) ,.ICEDI10 ( ICEDI10 ) ,.ICEDI9 ( ICEDI9 ) ,.ICEDI8 ( ICEDI8 )
 ,.ICEDI7 ( ICEDI7 ) ,.ICEDI6 ( ICEDI6 ) ,.ICEDI5 ( ICEDI5 ) ,.ICEDI4 ( ICEDI4 ) ,.ICEDI3 ( ICEDI3 ) ,.ICEDI2 ( ICEDI2 )
 ,.ICEDI1 ( ICEDI1 ) ,.ICEDI0 ( ICEDI0 ) ,.ICEWR ( ICEWR ) ,.ICERD ( ICERD ) ,.SYSRSOUTB ( SYSRSOUTB ) ,.SELEXMPC ( SELEXMPC )
 ,.SELRAMPC ( SELRAMPC ) ,.SELROMPC ( SELROMPC ) ,.SELBRAMPC ( SELBRAMPC ) ,.SELBFAPC ( SELBFAPC )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/mask.v
  MASK mask (
   .ICEDO31 ( ICEDOL31 ) ,.ICEDO23 ( ICEDOL23 ) ,.ICEDO15 ( ICEDOL15 ) ,.ICEDO30 ( ICEDOL30 ) ,.ICEDO22 ( ICEDOL22 ) ,.ICEDO14 ( ICEDOL14 ) ,.ICEDO29 ( ICEDOL29 )
 ,.ICEDO28 ( ICEDOL28 ) ,.ICEDO27 ( ICEDOL27 ) ,.ICEDO19 ( ICEDOL19 ) ,.ICEDO26 ( ICEDOL26 ) ,.ICEDO18 ( ICEDOL18 ) ,.ICEDO25 ( ICEDOL25 )
 ,.ICEDO17 ( ICEDOL17 ) ,.ICEDO24 ( ICEDOL24 ) ,.ICEDO16 ( ICEDOL16 ) ,.ICEDO21 ( ICEDOL21 ) ,.ICEDO13 ( ICEDOL13 ) ,.ICEDO20 ( ICEDOL20 )
 ,.ICEDO12 ( ICEDOL12 ) ,.ICEDO11 ( ICEDOL11 ) ,.ICEDO10 ( ICEDOL10 ) ,.ICEDO9 ( ICEDOL9 ) ,.ICEDO8 ( ICEDOL8 ) ,.ICEDO7 ( ICEDOL7 )
 ,.ICEDO6 ( ICEDOL6 ) ,.ICEDO5 ( ICEDOL5 ) ,.ICEDO4 ( ICEDOL4 ) ,.ICEDO3 ( ICEDOL3 ) ,.ICEDO2 ( ICEDOL2 ) ,.ICEDO1 ( ICEDOL1 )
 ,.ICEDO0 ( ICEDOL0 ) ,.SYSRSOUTB ( SYSRSOUTB ) ,.ICEIFA31 ( ICEIFA31 ) ,.ICEIFA23 ( ICEIFA23 ) ,.ICEIFA15 ( ICEIFA15 ) ,.ICEIFA30 ( ICEIFA30 )
 ,.ICEIFA22 ( ICEIFA22 ) ,.ICEIFA14 ( ICEIFA14 ) ,.ICEIFA29 ( ICEIFA29 ) ,.ICEIFA28 ( ICEIFA28 ) ,.ICEIFA27 ( ICEIFA27 ) ,.ICEIFA19 ( ICEIFA19 )
 ,.ICEIFA26 ( ICEIFA26 ) ,.ICEIFA18 ( ICEIFA18 ) ,.ICEIFA25 ( ICEIFA25 ) ,.ICEIFA17 ( ICEIFA17 ) ,.ICEIFA24 ( ICEIFA24 ) ,.ICEIFA16 ( ICEIFA16 )
 ,.ICEIFA21 ( ICEIFA21 ) ,.ICEIFA13 ( ICEIFA13 ) ,.ICEIFA20 ( ICEIFA20 ) ,.ICEIFA12 ( ICEIFA12 ) ,.ICEIFA11 ( ICEIFA11 ) ,.ICEIFA10 ( ICEIFA10 )
 ,.ICEIFA9 ( ICEIFA9 ) ,.ICEIFA8 ( ICEIFA8 ) ,.ICEIFA7 ( ICEIFA7 ) ,.ICEIFA6 ( ICEIFA6 ) ,.ICEIFA5 ( ICEIFA5 ) ,.ICEIFA4 ( ICEIFA4 )
 ,.ICEIFA3 ( ICEIFA3 ) ,.ICEIFA2 ( ICEIFA2 ) ,.ICEIFA1 ( ICEIFA1 ) ,.ICEIFA0 ( ICEIFA0 ) ,.ICEDI31 ( ICEDI31 ) ,.ICEDI23 ( ICEDI23 )
 ,.ICEDI15 ( ICEDI15 ) ,.ICEDI30 ( ICEDI30 ) ,.ICEDI22 ( ICEDI22 ) ,.ICEDI14 ( ICEDI14 ) ,.ICEDI29 ( ICEDI29 ) ,.ICEDI28 ( ICEDI28 )
 ,.ICEDI27 ( ICEDI27 ) ,.ICEDI19 ( ICEDI19 ) ,.ICEDI26 ( ICEDI26 ) ,.ICEDI18 ( ICEDI18 ) ,.ICEDI25 ( ICEDI25 ) ,.ICEDI17 ( ICEDI17 )
 ,.ICEDI24 ( ICEDI24 ) ,.ICEDI16 ( ICEDI16 ) ,.ICEDI21 ( ICEDI21 ) ,.ICEDI13 ( ICEDI13 ) ,.ICEDI20 ( ICEDI20 ) ,.ICEDI12 ( ICEDI12 )
 ,.ICEDI11 ( ICEDI11 ) ,.ICEDI10 ( ICEDI10 ) ,.ICEDI9 ( ICEDI9 ) ,.ICEDI8 ( ICEDI8 ) ,.ICEDI7 ( ICEDI7 ) ,.ICEDI6 ( ICEDI6 )
 ,.ICEDI5 ( ICEDI5 ) ,.ICEDI4 ( ICEDI4 ) ,.ICEDI3 ( ICEDI3 ) ,.ICEDI2 ( ICEDI2 ) ,.ICEDI1 ( ICEDI1 ) ,.ICEDI0 ( ICEDI0 )
 ,.ICEWR ( ICEWR ) ,.SVMODUSER ( SVMODUSER ) ,.ICEMSKRETRY ( ICEMSKRETRY ) ,.ICEMSKDBG ( ICEMSKDBG ) ,.ICEMSKWAIT ( ICEMSKWAIT ) ,.ICEMSKNMI ( ICEMSKNMI )
 ,.ICEMSKICE ( ICEMSKICE ) ,.ICEMSKTRAP ( ICEMSKTRAP ) ,.ICEMSKWDT ( ICEMSKWDT ) ,.ICEMSKLVI ( ICEMSKLVI ) ,.ICEMSKPOC ( ICEMSKPOC ) ,.ICEMSKTRST ( ICEMSKTRST )
 ,.ICEMSKTRSTFLG ( ICEMSKTRSTFLG )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/orbus-SS3rd.v
  ORBUS orbus (
   .MDR_RAM15 ( MDR_RAM15 ) ,.MDR_RAM14 ( MDR_RAM14 ) ,.MDR_RAM13 ( MDR_RAM13 ) ,.MDR_RAM12 ( MDR_RAM12 ) ,.MDR_RAM11 ( MDR_RAM11 ) ,.MDR_RAM10 ( MDR_RAM10 ) ,.MDR_RAM9 ( MDR_RAM9 )
 ,.MDR_RAM8 ( MDR_RAM8 ) ,.MDR_RAM7 ( MDR_RAM7 ) ,.MDR_RAM6 ( MDR_RAM6 ) ,.MDR_RAM5 ( MDR_RAM5 ) ,.MDR_RAM4 ( MDR_RAM4 ) ,.MDR_RAM3 ( MDR_RAM3 )
 ,.MDR_RAM2 ( MDR_RAM2 ) ,.MDR_RAM1 ( MDR_RAM1 ) ,.MDR_RAM0 ( MDR_RAM0 ) ,.MEMMDR15 ( MEMMDR15 ) ,.MEMMDR14 ( MEMMDR14 ) ,.MEMMDR13 ( MEMMDR13 )
 ,.MEMMDR12 ( MEMMDR12 ) ,.MEMMDR11 ( MEMMDR11 ) ,.MEMMDR10 ( MEMMDR10 ) ,.MEMMDR9 ( MEMMDR9 ) ,.MEMMDR8 ( MEMMDR8 ) ,.MEMMDR7 ( MEMMDR7 )
 ,.MEMMDR6 ( MEMMDR6 ) ,.MEMMDR5 ( MEMMDR5 ) ,.MEMMDR4 ( MEMMDR4 ) ,.MEMMDR3 ( MEMMDR3 ) ,.MEMMDR2 ( MEMMDR2 ) ,.MEMMDR1 ( MEMMDR1 )
 ,.MEMMDR0 ( MEMMDR0 ) ,.TRACEMDR15 ( TRACEMDR15 ) ,.TRACEMDR14 ( TRACEMDR14 ) ,.TRACEMDR13 ( TRACEMDR13 ) ,.TRACEMDR12 ( TRACEMDR12 ) ,.TRACEMDR11 ( TRACEMDR11 )
 ,.TRACEMDR10 ( TRACEMDR10 ) ,.TRACEMDR9 ( TRACEMDR9 ) ,.TRACEMDR8 ( TRACEMDR8 ) ,.TRACEMDR7 ( TRACEMDR7 ) ,.TRACEMDR6 ( TRACEMDR6 ) ,.TRACEMDR5 ( TRACEMDR5 )
 ,.TRACEMDR4 ( TRACEMDR4 ) ,.TRACEMDR3 ( TRACEMDR3 ) ,.TRACEMDR2 ( TRACEMDR2 ) ,.TRACEMDR1 ( TRACEMDR1 ) ,.TRACEMDR0 ( TRACEMDR0 ) ,.STATEMDR15 ( STATEMDR15 )
 ,.STATEMDR14 ( STATEMDR14 ) ,.STATEMDR13 ( STATEMDR13 ) ,.STATEMDR12 ( STATEMDR12 ) ,.STATEMDR11 ( STATEMDR11 ) ,.STATEMDR10 ( STATEMDR10 ) ,.STATEMDR9 ( STATEMDR9 )
 ,.STATEMDR8 ( STATEMDR8 ) ,.STATEMDR7 ( STATEMDR7 ) ,.STATEMDR6 ( STATEMDR6 ) ,.STATEMDR5 ( STATEMDR5 ) ,.STATEMDR4 ( STATEMDR4 ) ,.STATEMDR3 ( STATEMDR3 )
 ,.STATEMDR2 ( STATEMDR2 ) ,.STATEMDR1 ( STATEMDR1 ) ,.STATEMDR0 ( STATEMDR0 ) ,.BRKMDR15 ( BRKMDR15 ) ,.BRKMDR14 ( BRKMDR14 ) ,.BRKMDR13 ( BRKMDR13 )
 ,.BRKMDR12 ( BRKMDR12 ) ,.BRKMDR11 ( BRKMDR11 ) ,.BRKMDR10 ( BRKMDR10 ) ,.BRKMDR9 ( BRKMDR9 ) ,.BRKMDR8 ( BRKMDR8 ) ,.BRKMDR7 ( BRKMDR7 )
 ,.BRKMDR6 ( BRKMDR6 ) ,.BRKMDR5 ( BRKMDR5 ) ,.BRKMDR4 ( BRKMDR4 ) ,.BRKMDR3 ( BRKMDR3 ) ,.BRKMDR2 ( BRKMDR2 ) ,.BRKMDR1 ( BRKMDR1 )
 ,.BRKMDR0 ( BRKMDR0 ) ,.HOSTIFMDR15 ( HOSTIFMDR15 ) ,.HOSTIFMDR14 ( HOSTIFMDR14 ) ,.HOSTIFMDR13 ( HOSTIFMDR13 ) ,.HOSTIFMDR12 ( HOSTIFMDR12 ) ,.HOSTIFMDR11 ( HOSTIFMDR11 )
 ,.HOSTIFMDR10 ( HOSTIFMDR10 ) ,.HOSTIFMDR9 ( HOSTIFMDR9 ) ,.HOSTIFMDR8 ( HOSTIFMDR8 ) ,.HOSTIFMDR7 ( HOSTIFMDR7 ) ,.HOSTIFMDR6 ( HOSTIFMDR6 ) ,.HOSTIFMDR5 ( HOSTIFMDR5 )
 ,.HOSTIFMDR4 ( HOSTIFMDR4 ) ,.HOSTIFMDR3 ( HOSTIFMDR3 ) ,.HOSTIFMDR2 ( HOSTIFMDR2 ) ,.HOSTIFMDR1 ( HOSTIFMDR1 ) ,.HOSTIFMDR0 ( HOSTIFMDR0 ) ,.DFMDR15 ( DFMDR15 )
 ,.DFMDR14 ( DFMDR14 ) ,.DFMDR13 ( DFMDR13 ) ,.DFMDR12 ( DFMDR12 ) ,.DFMDR11 ( DFMDR11 ) ,.DFMDR10 ( DFMDR10 ) ,.DFMDR9 ( DFMDR9 )
 ,.DFMDR8 ( DFMDR8 ) ,.DFMDR7 ( DFMDR7 ) ,.DFMDR6 ( DFMDR6 ) ,.DFMDR5 ( DFMDR5 ) ,.DFMDR4 ( DFMDR4 ) ,.DFMDR3 ( DFMDR3 )
 ,.DFMDR2 ( DFMDR2 ) ,.DFMDR1 ( DFMDR1 ) ,.DFMDR0 ( DFMDR0 ) ,.SLDFLASH ( SLDFLASH )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/idversion.v
  IDVERSION idversion (
   .ICEDO31 ( ICEDOS31 ) ,.ICEDO23 ( ICEDOS23 ) ,.ICEDO15 ( ICEDOS15 ) ,.ICEDO30 ( ICEDOS30 ) ,.ICEDO22 ( ICEDOS22 ) ,.ICEDO14 ( ICEDOS14 ) ,.ICEDO29 ( ICEDOS29 )
 ,.ICEDO28 ( ICEDOS28 ) ,.ICEDO27 ( ICEDOS27 ) ,.ICEDO19 ( ICEDOS19 ) ,.ICEDO26 ( ICEDOS26 ) ,.ICEDO18 ( ICEDOS18 ) ,.ICEDO25 ( ICEDOS25 )
 ,.ICEDO17 ( ICEDOS17 ) ,.ICEDO24 ( ICEDOS24 ) ,.ICEDO16 ( ICEDOS16 ) ,.ICEDO21 ( ICEDOS21 ) ,.ICEDO13 ( ICEDOS13 ) ,.ICEDO20 ( ICEDOS20 )
 ,.ICEDO12 ( ICEDOS12 ) ,.ICEDO11 ( ICEDOS11 ) ,.ICEDO10 ( ICEDOS10 ) ,.ICEDO9 ( ICEDOS9 ) ,.ICEDO8 ( ICEDOS8 ) ,.ICEDO7 ( ICEDOS7 )
 ,.ICEDO6 ( ICEDOS6 ) ,.ICEDO5 ( ICEDOS5 ) ,.ICEDO4 ( ICEDOS4 ) ,.ICEDO3 ( ICEDOS3 ) ,.ICEDO2 ( ICEDOS2 ) ,.ICEDO1 ( ICEDOS1 )
 ,.ICEDO0 ( ICEDOS0 ) ,.IDVER31 ( IDVER31 ) ,.IDVER23 ( IDVER23 ) ,.IDVER15 ( IDVER15 ) ,.IDVER30 ( IDVER30 ) ,.IDVER22 ( IDVER22 )
 ,.IDVER14 ( IDVER14 ) ,.IDVER29 ( IDVER29 ) ,.IDVER28 ( IDVER28 ) ,.IDVER27 ( IDVER27 ) ,.IDVER19 ( IDVER19 ) ,.IDVER26 ( IDVER26 )
 ,.IDVER18 ( IDVER18 ) ,.IDVER25 ( IDVER25 ) ,.IDVER17 ( IDVER17 ) ,.IDVER24 ( IDVER24 ) ,.IDVER16 ( IDVER16 ) ,.IDVER21 ( IDVER21 )
 ,.IDVER13 ( IDVER13 ) ,.IDVER20 ( IDVER20 ) ,.IDVER12 ( IDVER12 ) ,.IDVER11 ( IDVER11 ) ,.IDVER10 ( IDVER10 ) ,.IDVER9 ( IDVER9 )
 ,.IDVER8 ( IDVER8 ) ,.IDVER7 ( IDVER7 ) ,.IDVER6 ( IDVER6 ) ,.IDVER5 ( IDVER5 ) ,.IDVER4 ( IDVER4 ) ,.IDVER3 ( IDVER3 )
 ,.IDVER2 ( IDVER2 ) ,.IDVER1 ( IDVER1 ) ,.IDVER0 ( IDVER0 ) ,.ICEIFA31 ( ICEIFA31 ) ,.ICEIFA23 ( ICEIFA23 ) ,.ICEIFA15 ( ICEIFA15 )
 ,.ICEIFA30 ( ICEIFA30 ) ,.ICEIFA22 ( ICEIFA22 ) ,.ICEIFA14 ( ICEIFA14 ) ,.ICEIFA29 ( ICEIFA29 ) ,.ICEIFA28 ( ICEIFA28 ) ,.ICEIFA27 ( ICEIFA27 )
 ,.ICEIFA19 ( ICEIFA19 ) ,.ICEIFA26 ( ICEIFA26 ) ,.ICEIFA18 ( ICEIFA18 ) ,.ICEIFA25 ( ICEIFA25 ) ,.ICEIFA17 ( ICEIFA17 ) ,.ICEIFA24 ( ICEIFA24 )
 ,.ICEIFA16 ( ICEIFA16 ) ,.ICEIFA21 ( ICEIFA21 ) ,.ICEIFA13 ( ICEIFA13 ) ,.ICEIFA20 ( ICEIFA20 ) ,.ICEIFA12 ( ICEIFA12 ) ,.ICEIFA11 ( ICEIFA11 )
 ,.ICEIFA10 ( ICEIFA10 ) ,.ICEIFA9 ( ICEIFA9 ) ,.ICEIFA8 ( ICEIFA8 ) ,.ICEIFA7 ( ICEIFA7 ) ,.ICEIFA6 ( ICEIFA6 ) ,.ICEIFA5 ( ICEIFA5 )
 ,.ICEIFA4 ( ICEIFA4 ) ,.ICEIFA3 ( ICEIFA3 ) ,.ICEIFA2 ( ICEIFA2 ) ,.ICEIFA1 ( ICEIFA1 ) ,.ICEIFA0 ( ICEIFA0 )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/test.v
  TESTCTL testctl (
   .ICEDO31 ( ICEDOT31 ) ,.ICEDO23 ( ICEDOT23 ) ,.ICEDO15 ( ICEDOT15 ) ,.ICEDO30 ( ICEDOT30 ) ,.ICEDO22 ( ICEDOT22 ) ,.ICEDO14 ( ICEDOT14 ) ,.ICEDO29 ( ICEDOT29 )
 ,.ICEDO28 ( ICEDOT28 ) ,.ICEDO27 ( ICEDOT27 ) ,.ICEDO19 ( ICEDOT19 ) ,.ICEDO26 ( ICEDOT26 ) ,.ICEDO18 ( ICEDOT18 ) ,.ICEDO25 ( ICEDOT25 )
 ,.ICEDO17 ( ICEDOT17 ) ,.ICEDO24 ( ICEDOT24 ) ,.ICEDO16 ( ICEDOT16 ) ,.ICEDO21 ( ICEDOT21 ) ,.ICEDO13 ( ICEDOT13 ) ,.ICEDO20 ( ICEDOT20 )
 ,.ICEDO12 ( ICEDOT12 ) ,.ICEDO11 ( ICEDOT11 ) ,.ICEDO10 ( ICEDOT10 ) ,.ICEDO9 ( ICEDOT9 ) ,.ICEDO8 ( ICEDOT8 ) ,.ICEDO7 ( ICEDOT7 )
 ,.ICEDO6 ( ICEDOT6 ) ,.ICEDO5 ( ICEDOT5 ) ,.ICEDO4 ( ICEDOT4 ) ,.ICEDO3 ( ICEDOT3 ) ,.ICEDO2 ( ICEDOT2 ) ,.ICEDO1 ( ICEDOT1 )
 ,.ICEDO0 ( ICEDOT0 ) ,.ICEIFA31 ( ICEIFA31 ) ,.ICEIFA23 ( ICEIFA23 ) ,.ICEIFA15 ( ICEIFA15 ) ,.ICEIFA30 ( ICEIFA30 ) ,.ICEIFA22 ( ICEIFA22 )
 ,.ICEIFA14 ( ICEIFA14 ) ,.ICEIFA29 ( ICEIFA29 ) ,.ICEIFA28 ( ICEIFA28 ) ,.ICEIFA27 ( ICEIFA27 ) ,.ICEIFA19 ( ICEIFA19 ) ,.ICEIFA26 ( ICEIFA26 )
 ,.ICEIFA18 ( ICEIFA18 ) ,.ICEIFA25 ( ICEIFA25 ) ,.ICEIFA17 ( ICEIFA17 ) ,.ICEIFA24 ( ICEIFA24 ) ,.ICEIFA16 ( ICEIFA16 ) ,.ICEIFA21 ( ICEIFA21 )
 ,.ICEIFA13 ( ICEIFA13 ) ,.ICEIFA20 ( ICEIFA20 ) ,.ICEIFA12 ( ICEIFA12 ) ,.ICEIFA11 ( ICEIFA11 ) ,.ICEIFA10 ( ICEIFA10 ) ,.ICEIFA9 ( ICEIFA9 )
 ,.ICEIFA8 ( ICEIFA8 ) ,.ICEIFA7 ( ICEIFA7 ) ,.ICEIFA6 ( ICEIFA6 ) ,.ICEIFA5 ( ICEIFA5 ) ,.ICEIFA4 ( ICEIFA4 ) ,.ICEIFA3 ( ICEIFA3 )
 ,.ICEIFA2 ( ICEIFA2 ) ,.ICEIFA1 ( ICEIFA1 ) ,.ICEIFA0 ( ICEIFA0 ) ,.ADDRTD144 ( ADDRTD144 ) ,.ADDRTD136 ( ADDRTD136 ) ,.ADDRTD128 ( ADDRTD128 )
 ,.ADDRTD143 ( ADDRTD143 ) ,.ADDRTD135 ( ADDRTD135 ) ,.ADDRTD127 ( ADDRTD127 ) ,.ADDRTD119 ( ADDRTD119 ) ,.ADDRTD142 ( ADDRTD142 ) ,.ADDRTD134 ( ADDRTD134 )
 ,.ADDRTD126 ( ADDRTD126 ) ,.ADDRTD118 ( ADDRTD118 ) ,.ADDRTD141 ( ADDRTD141 ) ,.ADDRTD133 ( ADDRTD133 ) ,.ADDRTD125 ( ADDRTD125 ) ,.ADDRTD117 ( ADDRTD117 )
 ,.ADDRTD109 ( ADDRTD109 ) ,.ADDRTD140 ( ADDRTD140 ) ,.ADDRTD132 ( ADDRTD132 ) ,.ADDRTD124 ( ADDRTD124 ) ,.ADDRTD116 ( ADDRTD116 ) ,.ADDRTD108 ( ADDRTD108 )
 ,.ADDRTD139 ( ADDRTD139 ) ,.ADDRTD138 ( ADDRTD138 ) ,.ADDRTD137 ( ADDRTD137 ) ,.ADDRTD129 ( ADDRTD129 ) ,.ADDRTD131 ( ADDRTD131 ) ,.ADDRTD123 ( ADDRTD123 )
 ,.ADDRTD115 ( ADDRTD115 ) ,.ADDRTD107 ( ADDRTD107 ) ,.ADDRTD130 ( ADDRTD130 ) ,.ADDRTD122 ( ADDRTD122 ) ,.ADDRTD114 ( ADDRTD114 ) ,.ADDRTD106 ( ADDRTD106 )
 ,.ADDRTD121 ( ADDRTD121 ) ,.ADDRTD113 ( ADDRTD113 ) ,.ADDRTD105 ( ADDRTD105 ) ,.ADDRTD120 ( ADDRTD120 ) ,.ADDRTD112 ( ADDRTD112 ) ,.ADDRTD104 ( ADDRTD104 )
 ,.ADDRTD111 ( ADDRTD111 ) ,.ADDRTD103 ( ADDRTD103 ) ,.ADDRTD110 ( ADDRTD110 ) ,.ADDRTD102 ( ADDRTD102 ) ,.ADDRTD101 ( ADDRTD101 ) ,.ADDRTD100 ( ADDRTD100 )
 ,.ADDRTD99 ( ADDRTD99 ) ,.ADDRTD98 ( ADDRTD98 ) ,.ADDRTD97 ( ADDRTD97 ) ,.ADDRTD89 ( ADDRTD89 ) ,.ADDRTD96 ( ADDRTD96 ) ,.ADDRTD88 ( ADDRTD88 )
 ,.ADDRTD95 ( ADDRTD95 ) ,.ADDRTD87 ( ADDRTD87 ) ,.ADDRTD79 ( ADDRTD79 ) ,.ADDRTD94 ( ADDRTD94 ) ,.ADDRTD86 ( ADDRTD86 ) ,.ADDRTD78 ( ADDRTD78 )
 ,.ADDRTD93 ( ADDRTD93 ) ,.ADDRTD85 ( ADDRTD85 ) ,.ADDRTD77 ( ADDRTD77 ) ,.ADDRTD69 ( ADDRTD69 ) ,.ADDRTD92 ( ADDRTD92 ) ,.ADDRTD84 ( ADDRTD84 )
 ,.ADDRTD76 ( ADDRTD76 ) ,.ADDRTD68 ( ADDRTD68 ) ,.ADDRTD91 ( ADDRTD91 ) ,.ADDRTD83 ( ADDRTD83 ) ,.ADDRTD75 ( ADDRTD75 ) ,.ADDRTD67 ( ADDRTD67 )
 ,.ADDRTD59 ( ADDRTD59 ) ,.ADDRTD90 ( ADDRTD90 ) ,.ADDRTD82 ( ADDRTD82 ) ,.ADDRTD74 ( ADDRTD74 ) ,.ADDRTD66 ( ADDRTD66 ) ,.ADDRTD58 ( ADDRTD58 )
 ,.ADDRTD81 ( ADDRTD81 ) ,.ADDRTD73 ( ADDRTD73 ) ,.ADDRTD65 ( ADDRTD65 ) ,.ADDRTD57 ( ADDRTD57 ) ,.ADDRTD49 ( ADDRTD49 ) ,.ADDRTD80 ( ADDRTD80 )
 ,.ADDRTD72 ( ADDRTD72 ) ,.ADDRTD64 ( ADDRTD64 ) ,.ADDRTD56 ( ADDRTD56 ) ,.ADDRTD48 ( ADDRTD48 ) ,.ADDRTD71 ( ADDRTD71 ) ,.ADDRTD63 ( ADDRTD63 )
 ,.ADDRTD55 ( ADDRTD55 ) ,.ADDRTD47 ( ADDRTD47 ) ,.ADDRTD39 ( ADDRTD39 ) ,.ADDRTD70 ( ADDRTD70 ) ,.ADDRTD62 ( ADDRTD62 ) ,.ADDRTD54 ( ADDRTD54 )
 ,.ADDRTD46 ( ADDRTD46 ) ,.ADDRTD38 ( ADDRTD38 ) ,.ADDRTD61 ( ADDRTD61 ) ,.ADDRTD53 ( ADDRTD53 ) ,.ADDRTD45 ( ADDRTD45 ) ,.ADDRTD37 ( ADDRTD37 )
 ,.ADDRTD29 ( ADDRTD29 ) ,.ADDRTD60 ( ADDRTD60 ) ,.ADDRTD52 ( ADDRTD52 ) ,.ADDRTD44 ( ADDRTD44 ) ,.ADDRTD36 ( ADDRTD36 ) ,.ADDRTD28 ( ADDRTD28 )
 ,.ADDRTD51 ( ADDRTD51 ) ,.ADDRTD43 ( ADDRTD43 ) ,.ADDRTD35 ( ADDRTD35 ) ,.ADDRTD27 ( ADDRTD27 ) ,.ADDRTD19 ( ADDRTD19 ) ,.ADDRTD50 ( ADDRTD50 )
 ,.ADDRTD42 ( ADDRTD42 ) ,.ADDRTD34 ( ADDRTD34 ) ,.ADDRTD26 ( ADDRTD26 ) ,.ADDRTD18 ( ADDRTD18 ) ,.ADDRTD41 ( ADDRTD41 ) ,.ADDRTD33 ( ADDRTD33 )
 ,.ADDRTD25 ( ADDRTD25 ) ,.ADDRTD17 ( ADDRTD17 ) ,.ADDRTD40 ( ADDRTD40 ) ,.ADDRTD32 ( ADDRTD32 ) ,.ADDRTD24 ( ADDRTD24 ) ,.ADDRTD16 ( ADDRTD16 )
 ,.ADDRTD31 ( ADDRTD31 ) ,.ADDRTD23 ( ADDRTD23 ) ,.ADDRTD15 ( ADDRTD15 ) ,.ADDRTD30 ( ADDRTD30 ) ,.ADDRTD22 ( ADDRTD22 ) ,.ADDRTD14 ( ADDRTD14 )
 ,.ADDRTD21 ( ADDRTD21 ) ,.ADDRTD13 ( ADDRTD13 ) ,.ADDRTD20 ( ADDRTD20 ) ,.ADDRTD12 ( ADDRTD12 ) ,.ADDRTD11 ( ADDRTD11 ) ,.ADDRTD10 ( ADDRTD10 )
 ,.ADDRTD9 ( ADDRTD9 ) ,.ADDRTD8 ( ADDRTD8 ) ,.ADDRTD7 ( ADDRTD7 ) ,.ADDRTD6 ( ADDRTD6 ) ,.ADDRTD5 ( ADDRTD5 ) ,.ADDRTD4 ( ADDRTD4 )
 ,.ADDRTD3 ( ADDRTD3 ) ,.ADDRTD2 ( ADDRTD2 ) ,.ADDRTD1 ( ADDRTD1 ) ,.ADDRICE11 ( ADDRICE11 ) ,.ADDRICE10 ( ADDRICE10 ) ,.ADDRICE9 ( ADDRICE9 )
 ,.ADDRICE8 ( ADDRICE8 ) ,.ADDRICE7 ( ADDRICE7 ) ,.ADDRICE6 ( ADDRICE6 ) ,.ADDRICE5 ( ADDRICE5 ) ,.ADDRICE4 ( ADDRICE4 ) ,.ADDRICE3 ( ADDRICE3 )
 ,.ADDRICE2 ( ADDRICE2 ) ,.ADDRICE1 ( ADDRICE1 ) ,.ADDRICE0 ( ADDRICE0 ) ,.ADDRPINRD ( ADDRPINRD ) ,.ADDRPINMD ( ADDRPINMD ) ,.ADDRPINLV ( ADDRPINLV )
 ,.TP144D3 ( TP144D3 ) ,.TP136D3 ( TP136D3 ) ,.TP128D3 ( TP128D3 ) ,.TP144D2 ( TP144D2 ) ,.TP136D2 ( TP136D2 ) ,.TP128D2 ( TP128D2 )
 ,.TP144D1 ( TP144D1 ) ,.TP136D1 ( TP136D1 ) ,.TP128D1 ( TP128D1 ) ,.TP144D0 ( TP144D0 ) ,.TP136D0 ( TP136D0 ) ,.TP128D0 ( TP128D0 )
 ,.TP143D3 ( TP143D3 ) ,.TP135D3 ( TP135D3 ) ,.TP127D3 ( TP127D3 ) ,.TP119D3 ( TP119D3 ) ,.TP143D2 ( TP143D2 ) ,.TP135D2 ( TP135D2 )
 ,.TP127D2 ( TP127D2 ) ,.TP119D2 ( TP119D2 ) ,.TP143D1 ( TP143D1 ) ,.TP135D1 ( TP135D1 ) ,.TP127D1 ( TP127D1 ) ,.TP119D1 ( TP119D1 )
 ,.TP143D0 ( TP143D0 ) ,.TP135D0 ( TP135D0 ) ,.TP127D0 ( TP127D0 ) ,.TP119D0 ( TP119D0 ) ,.TP142D3 ( TP142D3 ) ,.TP134D3 ( TP134D3 )
 ,.TP126D3 ( TP126D3 ) ,.TP118D3 ( TP118D3 ) ,.TP142D2 ( TP142D2 ) ,.TP134D2 ( TP134D2 ) ,.TP126D2 ( TP126D2 ) ,.TP118D2 ( TP118D2 )
 ,.TP142D1 ( TP142D1 ) ,.TP134D1 ( TP134D1 ) ,.TP126D1 ( TP126D1 ) ,.TP118D1 ( TP118D1 ) ,.TP142D0 ( TP142D0 ) ,.TP134D0 ( TP134D0 )
 ,.TP126D0 ( TP126D0 ) ,.TP118D0 ( TP118D0 ) ,.TP141D3 ( TP141D3 ) ,.TP133D3 ( TP133D3 ) ,.TP125D3 ( TP125D3 ) ,.TP117D3 ( TP117D3 )
 ,.TP109D3 ( TP109D3 ) ,.TP141D2 ( TP141D2 ) ,.TP133D2 ( TP133D2 ) ,.TP125D2 ( TP125D2 ) ,.TP117D2 ( TP117D2 ) ,.TP109D2 ( TP109D2 )
 ,.TP141D1 ( TP141D1 ) ,.TP133D1 ( TP133D1 ) ,.TP125D1 ( TP125D1 ) ,.TP117D1 ( TP117D1 ) ,.TP109D1 ( TP109D1 ) ,.TP141D0 ( TP141D0 )
 ,.TP133D0 ( TP133D0 ) ,.TP125D0 ( TP125D0 ) ,.TP117D0 ( TP117D0 ) ,.TP109D0 ( TP109D0 ) ,.TP140D3 ( TP140D3 ) ,.TP132D3 ( TP132D3 )
 ,.TP124D3 ( TP124D3 ) ,.TP116D3 ( TP116D3 ) ,.TP108D3 ( TP108D3 ) ,.TP140D2 ( TP140D2 ) ,.TP132D2 ( TP132D2 ) ,.TP124D2 ( TP124D2 )
 ,.TP116D2 ( TP116D2 ) ,.TP108D2 ( TP108D2 ) ,.TP140D1 ( TP140D1 ) ,.TP132D1 ( TP132D1 ) ,.TP124D1 ( TP124D1 ) ,.TP116D1 ( TP116D1 )
 ,.TP108D1 ( TP108D1 ) ,.TP140D0 ( TP140D0 ) ,.TP132D0 ( TP132D0 ) ,.TP124D0 ( TP124D0 ) ,.TP116D0 ( TP116D0 ) ,.TP108D0 ( TP108D0 )
 ,.TP139D3 ( TP139D3 ) ,.TP139D2 ( TP139D2 ) ,.TP139D1 ( TP139D1 ) ,.TP139D0 ( TP139D0 ) ,.TP138D3 ( TP138D3 ) ,.TP138D2 ( TP138D2 )
 ,.TP138D1 ( TP138D1 ) ,.TP138D0 ( TP138D0 ) ,.TP137D3 ( TP137D3 ) ,.TP129D3 ( TP129D3 ) ,.TP137D2 ( TP137D2 ) ,.TP129D2 ( TP129D2 )
 ,.TP137D1 ( TP137D1 ) ,.TP129D1 ( TP129D1 ) ,.TP137D0 ( TP137D0 ) ,.TP129D0 ( TP129D0 ) ,.TP131D3 ( TP131D3 ) ,.TP123D3 ( TP123D3 )
 ,.TP115D3 ( TP115D3 ) ,.TP107D3 ( TP107D3 ) ,.TP131D2 ( TP131D2 ) ,.TP123D2 ( TP123D2 ) ,.TP115D2 ( TP115D2 ) ,.TP107D2 ( TP107D2 )
 ,.TP131D1 ( TP131D1 ) ,.TP123D1 ( TP123D1 ) ,.TP115D1 ( TP115D1 ) ,.TP107D1 ( TP107D1 ) ,.TP131D0 ( TP131D0 ) ,.TP123D0 ( TP123D0 )
 ,.TP115D0 ( TP115D0 ) ,.TP107D0 ( TP107D0 ) ,.TP130D3 ( TP130D3 ) ,.TP122D3 ( TP122D3 ) ,.TP114D3 ( TP114D3 ) ,.TP106D3 ( TP106D3 )
 ,.TP130D2 ( TP130D2 ) ,.TP122D2 ( TP122D2 ) ,.TP114D2 ( TP114D2 ) ,.TP106D2 ( TP106D2 ) ,.TP130D1 ( TP130D1 ) ,.TP122D1 ( TP122D1 )
 ,.TP114D1 ( TP114D1 ) ,.TP106D1 ( TP106D1 ) ,.TP130D0 ( TP130D0 ) ,.TP122D0 ( TP122D0 ) ,.TP114D0 ( TP114D0 ) ,.TP106D0 ( TP106D0 )
 ,.TP121D3 ( TP121D3 ) ,.TP113D3 ( TP113D3 ) ,.TP105D3 ( TP105D3 ) ,.TP121D2 ( TP121D2 ) ,.TP113D2 ( TP113D2 ) ,.TP105D2 ( TP105D2 )
 ,.TP121D1 ( TP121D1 ) ,.TP113D1 ( TP113D1 ) ,.TP105D1 ( TP105D1 ) ,.TP121D0 ( TP121D0 ) ,.TP113D0 ( TP113D0 ) ,.TP105D0 ( TP105D0 )
 ,.TP120D3 ( TP120D3 ) ,.TP112D3 ( TP112D3 ) ,.TP104D3 ( TP104D3 ) ,.TP120D2 ( TP120D2 ) ,.TP112D2 ( TP112D2 ) ,.TP104D2 ( TP104D2 )
 ,.TP120D1 ( TP120D1 ) ,.TP112D1 ( TP112D1 ) ,.TP104D1 ( TP104D1 ) ,.TP120D0 ( TP120D0 ) ,.TP112D0 ( TP112D0 ) ,.TP104D0 ( TP104D0 )
 ,.TP111D3 ( TP111D3 ) ,.TP103D3 ( TP103D3 ) ,.TP111D2 ( TP111D2 ) ,.TP103D2 ( TP103D2 ) ,.TP111D1 ( TP111D1 ) ,.TP103D1 ( TP103D1 )
 ,.TP111D0 ( TP111D0 ) ,.TP103D0 ( TP103D0 ) ,.TP110D3 ( TP110D3 ) ,.TP102D3 ( TP102D3 ) ,.TP110D2 ( TP110D2 ) ,.TP102D2 ( TP102D2 )
 ,.TP110D1 ( TP110D1 ) ,.TP102D1 ( TP102D1 ) ,.TP110D0 ( TP110D0 ) ,.TP102D0 ( TP102D0 ) ,.TP101D3 ( TP101D3 ) ,.TP101D2 ( TP101D2 )
 ,.TP101D1 ( TP101D1 ) ,.TP101D0 ( TP101D0 ) ,.TP100D3 ( TP100D3 ) ,.TP100D2 ( TP100D2 ) ,.TP100D1 ( TP100D1 ) ,.TP100D0 ( TP100D0 )
 ,.TP99D3 ( TP99D3 ) ,.TP99D2 ( TP99D2 ) ,.TP99D1 ( TP99D1 ) ,.TP99D0 ( TP99D0 ) ,.TP98D3 ( TP98D3 ) ,.TP98D2 ( TP98D2 )
 ,.TP98D1 ( TP98D1 ) ,.TP98D0 ( TP98D0 ) ,.TP97D3 ( TP97D3 ) ,.TP89D3 ( TP89D3 ) ,.TP97D2 ( TP97D2 ) ,.TP89D2 ( TP89D2 )
 ,.TP97D1 ( TP97D1 ) ,.TP89D1 ( TP89D1 ) ,.TP97D0 ( TP97D0 ) ,.TP89D0 ( TP89D0 ) ,.TP96D3 ( TP96D3 ) ,.TP88D3 ( TP88D3 )
 ,.TP96D2 ( TP96D2 ) ,.TP88D2 ( TP88D2 ) ,.TP96D1 ( TP96D1 ) ,.TP88D1 ( TP88D1 ) ,.TP96D0 ( TP96D0 ) ,.TP88D0 ( TP88D0 )
 ,.TP95D3 ( TP95D3 ) ,.TP87D3 ( TP87D3 ) ,.TP79D3 ( TP79D3 ) ,.TP95D2 ( TP95D2 ) ,.TP87D2 ( TP87D2 ) ,.TP79D2 ( TP79D2 )
 ,.TP95D1 ( TP95D1 ) ,.TP87D1 ( TP87D1 ) ,.TP79D1 ( TP79D1 ) ,.TP95D0 ( TP95D0 ) ,.TP87D0 ( TP87D0 ) ,.TP79D0 ( TP79D0 )
 ,.TP94D3 ( TP94D3 ) ,.TP86D3 ( TP86D3 ) ,.TP78D3 ( TP78D3 ) ,.TP94D2 ( TP94D2 ) ,.TP86D2 ( TP86D2 ) ,.TP78D2 ( TP78D2 )
 ,.TP94D1 ( TP94D1 ) ,.TP86D1 ( TP86D1 ) ,.TP78D1 ( TP78D1 ) ,.TP94D0 ( TP94D0 ) ,.TP86D0 ( TP86D0 ) ,.TP78D0 ( TP78D0 )
 ,.TP93D3 ( TP93D3 ) ,.TP85D3 ( TP85D3 ) ,.TP77D3 ( TP77D3 ) ,.TP69D3 ( TP69D3 ) ,.TP93D2 ( TP93D2 ) ,.TP85D2 ( TP85D2 )
 ,.TP77D2 ( TP77D2 ) ,.TP69D2 ( TP69D2 ) ,.TP93D1 ( TP93D1 ) ,.TP85D1 ( TP85D1 ) ,.TP77D1 ( TP77D1 ) ,.TP69D1 ( TP69D1 )
 ,.TP93D0 ( TP93D0 ) ,.TP85D0 ( TP85D0 ) ,.TP77D0 ( TP77D0 ) ,.TP69D0 ( TP69D0 ) ,.TP92D3 ( TP92D3 ) ,.TP84D3 ( TP84D3 )
 ,.TP76D3 ( TP76D3 ) ,.TP68D3 ( TP68D3 ) ,.TP92D2 ( TP92D2 ) ,.TP84D2 ( TP84D2 ) ,.TP76D2 ( TP76D2 ) ,.TP68D2 ( TP68D2 )
 ,.TP92D1 ( TP92D1 ) ,.TP84D1 ( TP84D1 ) ,.TP76D1 ( TP76D1 ) ,.TP68D1 ( TP68D1 ) ,.TP92D0 ( TP92D0 ) ,.TP84D0 ( TP84D0 )
 ,.TP76D0 ( TP76D0 ) ,.TP68D0 ( TP68D0 ) ,.TP91D3 ( TP91D3 ) ,.TP83D3 ( TP83D3 ) ,.TP75D3 ( TP75D3 ) ,.TP67D3 ( TP67D3 )
 ,.TP59D3 ( TP59D3 ) ,.TP91D2 ( TP91D2 ) ,.TP83D2 ( TP83D2 ) ,.TP75D2 ( TP75D2 ) ,.TP67D2 ( TP67D2 ) ,.TP59D2 ( TP59D2 )
 ,.TP91D1 ( TP91D1 ) ,.TP83D1 ( TP83D1 ) ,.TP75D1 ( TP75D1 ) ,.TP67D1 ( TP67D1 ) ,.TP59D1 ( TP59D1 ) ,.TP91D0 ( TP91D0 )
 ,.TP83D0 ( TP83D0 ) ,.TP75D0 ( TP75D0 ) ,.TP67D0 ( TP67D0 ) ,.TP59D0 ( TP59D0 ) ,.TP90D3 ( TP90D3 ) ,.TP82D3 ( TP82D3 )
 ,.TP74D3 ( TP74D3 ) ,.TP66D3 ( TP66D3 ) ,.TP58D3 ( TP58D3 ) ,.TP90D2 ( TP90D2 ) ,.TP82D2 ( TP82D2 ) ,.TP74D2 ( TP74D2 )
 ,.TP66D2 ( TP66D2 ) ,.TP58D2 ( TP58D2 ) ,.TP90D1 ( TP90D1 ) ,.TP82D1 ( TP82D1 ) ,.TP74D1 ( TP74D1 ) ,.TP66D1 ( TP66D1 )
 ,.TP58D1 ( TP58D1 ) ,.TP90D0 ( TP90D0 ) ,.TP82D0 ( TP82D0 ) ,.TP74D0 ( TP74D0 ) ,.TP66D0 ( TP66D0 ) ,.TP58D0 ( TP58D0 )
 ,.TP81D3 ( TP81D3 ) ,.TP73D3 ( TP73D3 ) ,.TP65D3 ( TP65D3 ) ,.TP57D3 ( TP57D3 ) ,.TP49D3 ( TP49D3 ) ,.TP81D2 ( TP81D2 )
 ,.TP73D2 ( TP73D2 ) ,.TP65D2 ( TP65D2 ) ,.TP57D2 ( TP57D2 ) ,.TP49D2 ( TP49D2 ) ,.TP81D1 ( TP81D1 ) ,.TP73D1 ( TP73D1 )
 ,.TP65D1 ( TP65D1 ) ,.TP57D1 ( TP57D1 ) ,.TP49D1 ( TP49D1 ) ,.TP81D0 ( TP81D0 ) ,.TP73D0 ( TP73D0 ) ,.TP65D0 ( TP65D0 )
 ,.TP57D0 ( TP57D0 ) ,.TP49D0 ( TP49D0 ) ,.TP80D3 ( TP80D3 ) ,.TP72D3 ( TP72D3 ) ,.TP64D3 ( TP64D3 ) ,.TP56D3 ( TP56D3 )
 ,.TP48D3 ( TP48D3 ) ,.TP80D2 ( TP80D2 ) ,.TP72D2 ( TP72D2 ) ,.TP64D2 ( TP64D2 ) ,.TP56D2 ( TP56D2 ) ,.TP48D2 ( TP48D2 )
 ,.TP80D1 ( TP80D1 ) ,.TP72D1 ( TP72D1 ) ,.TP64D1 ( TP64D1 ) ,.TP56D1 ( TP56D1 ) ,.TP48D1 ( TP48D1 ) ,.TP80D0 ( TP80D0 )
 ,.TP72D0 ( TP72D0 ) ,.TP64D0 ( TP64D0 ) ,.TP56D0 ( TP56D0 ) ,.TP48D0 ( TP48D0 ) ,.TP71D3 ( TP71D3 ) ,.TP63D3 ( TP63D3 )
 ,.TP55D3 ( TP55D3 ) ,.TP47D3 ( TP47D3 ) ,.TP39D3 ( TP39D3 ) ,.TP71D2 ( TP71D2 ) ,.TP63D2 ( TP63D2 ) ,.TP55D2 ( TP55D2 )
 ,.TP47D2 ( TP47D2 ) ,.TP39D2 ( TP39D2 ) ,.TP71D1 ( TP71D1 ) ,.TP63D1 ( TP63D1 ) ,.TP55D1 ( TP55D1 ) ,.TP47D1 ( TP47D1 )
 ,.TP39D1 ( TP39D1 ) ,.TP71D0 ( TP71D0 ) ,.TP63D0 ( TP63D0 ) ,.TP55D0 ( TP55D0 ) ,.TP47D0 ( TP47D0 ) ,.TP39D0 ( TP39D0 )
 ,.TP70D3 ( TP70D3 ) ,.TP62D3 ( TP62D3 ) ,.TP54D3 ( TP54D3 ) ,.TP46D3 ( TP46D3 ) ,.TP38D3 ( TP38D3 ) ,.TP70D2 ( TP70D2 )
 ,.TP62D2 ( TP62D2 ) ,.TP54D2 ( TP54D2 ) ,.TP46D2 ( TP46D2 ) ,.TP38D2 ( TP38D2 ) ,.TP70D1 ( TP70D1 ) ,.TP62D1 ( TP62D1 )
 ,.TP54D1 ( TP54D1 ) ,.TP46D1 ( TP46D1 ) ,.TP38D1 ( TP38D1 ) ,.TP70D0 ( TP70D0 ) ,.TP62D0 ( TP62D0 ) ,.TP54D0 ( TP54D0 )
 ,.TP46D0 ( TP46D0 ) ,.TP38D0 ( TP38D0 ) ,.TP61D3 ( TP61D3 ) ,.TP53D3 ( TP53D3 ) ,.TP45D3 ( TP45D3 ) ,.TP37D3 ( TP37D3 )
 ,.TP29D3 ( TP29D3 ) ,.TP61D2 ( TP61D2 ) ,.TP53D2 ( TP53D2 ) ,.TP45D2 ( TP45D2 ) ,.TP37D2 ( TP37D2 ) ,.TP29D2 ( TP29D2 )
 ,.TP61D1 ( TP61D1 ) ,.TP53D1 ( TP53D1 ) ,.TP45D1 ( TP45D1 ) ,.TP37D1 ( TP37D1 ) ,.TP29D1 ( TP29D1 ) ,.TP61D0 ( TP61D0 )
 ,.TP53D0 ( TP53D0 ) ,.TP45D0 ( TP45D0 ) ,.TP37D0 ( TP37D0 ) ,.TP29D0 ( TP29D0 ) ,.TP60D3 ( TP60D3 ) ,.TP52D3 ( TP52D3 )
 ,.TP44D3 ( TP44D3 ) ,.TP36D3 ( TP36D3 ) ,.TP28D3 ( TP28D3 ) ,.TP60D2 ( TP60D2 ) ,.TP52D2 ( TP52D2 ) ,.TP44D2 ( TP44D2 )
 ,.TP36D2 ( TP36D2 ) ,.TP28D2 ( TP28D2 ) ,.TP60D1 ( TP60D1 ) ,.TP52D1 ( TP52D1 ) ,.TP44D1 ( TP44D1 ) ,.TP36D1 ( TP36D1 )
 ,.TP28D1 ( TP28D1 ) ,.TP60D0 ( TP60D0 ) ,.TP52D0 ( TP52D0 ) ,.TP44D0 ( TP44D0 ) ,.TP36D0 ( TP36D0 ) ,.TP28D0 ( TP28D0 )
 ,.TP51D3 ( TP51D3 ) ,.TP43D3 ( TP43D3 ) ,.TP35D3 ( TP35D3 ) ,.TP27D3 ( TP27D3 ) ,.TP19D3 ( TP19D3 ) ,.TP51D2 ( TP51D2 )
 ,.TP43D2 ( TP43D2 ) ,.TP35D2 ( TP35D2 ) ,.TP27D2 ( TP27D2 ) ,.TP19D2 ( TP19D2 ) ,.TP51D1 ( TP51D1 ) ,.TP43D1 ( TP43D1 )
 ,.TP35D1 ( TP35D1 ) ,.TP27D1 ( TP27D1 ) ,.TP19D1 ( TP19D1 ) ,.TP51D0 ( TP51D0 ) ,.TP43D0 ( TP43D0 ) ,.TP35D0 ( TP35D0 )
 ,.TP27D0 ( TP27D0 ) ,.TP19D0 ( TP19D0 ) ,.TP50D3 ( TP50D3 ) ,.TP42D3 ( TP42D3 ) ,.TP34D3 ( TP34D3 ) ,.TP26D3 ( TP26D3 )
 ,.TP18D3 ( TP18D3 ) ,.TP50D2 ( TP50D2 ) ,.TP42D2 ( TP42D2 ) ,.TP34D2 ( TP34D2 ) ,.TP26D2 ( TP26D2 ) ,.TP18D2 ( TP18D2 )
 ,.TP50D1 ( TP50D1 ) ,.TP42D1 ( TP42D1 ) ,.TP34D1 ( TP34D1 ) ,.TP26D1 ( TP26D1 ) ,.TP18D1 ( TP18D1 ) ,.TP50D0 ( TP50D0 )
 ,.TP42D0 ( TP42D0 ) ,.TP34D0 ( TP34D0 ) ,.TP26D0 ( TP26D0 ) ,.TP18D0 ( TP18D0 ) ,.TP41D3 ( TP41D3 ) ,.TP33D3 ( TP33D3 )
 ,.TP25D3 ( TP25D3 ) ,.TP17D3 ( TP17D3 ) ,.TP41D2 ( TP41D2 ) ,.TP33D2 ( TP33D2 ) ,.TP25D2 ( TP25D2 ) ,.TP17D2 ( TP17D2 )
 ,.TP41D1 ( TP41D1 ) ,.TP33D1 ( TP33D1 ) ,.TP25D1 ( TP25D1 ) ,.TP17D1 ( TP17D1 ) ,.TP41D0 ( TP41D0 ) ,.TP33D0 ( TP33D0 )
 ,.TP25D0 ( TP25D0 ) ,.TP17D0 ( TP17D0 ) ,.TP40D3 ( TP40D3 ) ,.TP32D3 ( TP32D3 ) ,.TP24D3 ( TP24D3 ) ,.TP16D3 ( TP16D3 )
 ,.TP40D2 ( TP40D2 ) ,.TP32D2 ( TP32D2 ) ,.TP24D2 ( TP24D2 ) ,.TP16D2 ( TP16D2 ) ,.TP40D1 ( TP40D1 ) ,.TP32D1 ( TP32D1 )
 ,.TP24D1 ( TP24D1 ) ,.TP16D1 ( TP16D1 ) ,.TP40D0 ( TP40D0 ) ,.TP32D0 ( TP32D0 ) ,.TP24D0 ( TP24D0 ) ,.TP16D0 ( TP16D0 )
 ,.TP31D3 ( TP31D3 ) ,.TP23D3 ( TP23D3 ) ,.TP15D3 ( TP15D3 ) ,.TP31D2 ( TP31D2 ) ,.TP23D2 ( TP23D2 ) ,.TP15D2 ( TP15D2 )
 ,.TP31D1 ( TP31D1 ) ,.TP23D1 ( TP23D1 ) ,.TP15D1 ( TP15D1 ) ,.TP31D0 ( TP31D0 ) ,.TP23D0 ( TP23D0 ) ,.TP15D0 ( TP15D0 )
 ,.TP30D3 ( TP30D3 ) ,.TP22D3 ( TP22D3 ) ,.TP14D3 ( TP14D3 ) ,.TP30D2 ( TP30D2 ) ,.TP22D2 ( TP22D2 ) ,.TP14D2 ( TP14D2 )
 ,.TP30D1 ( TP30D1 ) ,.TP22D1 ( TP22D1 ) ,.TP14D1 ( TP14D1 ) ,.TP30D0 ( TP30D0 ) ,.TP22D0 ( TP22D0 ) ,.TP14D0 ( TP14D0 )
 ,.TP21D3 ( TP21D3 ) ,.TP13D3 ( TP13D3 ) ,.TP21D2 ( TP21D2 ) ,.TP13D2 ( TP13D2 ) ,.TP21D1 ( TP21D1 ) ,.TP13D1 ( TP13D1 )
 ,.TP21D0 ( TP21D0 ) ,.TP13D0 ( TP13D0 ) ,.TP20D3 ( TP20D3 ) ,.TP12D3 ( TP12D3 ) ,.TP20D2 ( TP20D2 ) ,.TP12D2 ( TP12D2 )
 ,.TP20D1 ( TP20D1 ) ,.TP12D1 ( TP12D1 ) ,.TP20D0 ( TP20D0 ) ,.TP12D0 ( TP12D0 ) ,.TP11D3 ( TP11D3 ) ,.TP11D2 ( TP11D2 )
 ,.TP11D1 ( TP11D1 ) ,.TP11D0 ( TP11D0 ) ,.TP10D3 ( TP10D3 ) ,.TP10D2 ( TP10D2 ) ,.TP10D1 ( TP10D1 ) ,.TP10D0 ( TP10D0 )
 ,.TP9D3 ( TP9D3 ) ,.TP9D2 ( TP9D2 ) ,.TP9D1 ( TP9D1 ) ,.TP9D0 ( TP9D0 ) ,.TP8D3 ( TP8D3 ) ,.TP8D2 ( TP8D2 )
 ,.TP8D1 ( TP8D1 ) ,.TP8D0 ( TP8D0 ) ,.TP7D3 ( TP7D3 ) ,.TP7D2 ( TP7D2 ) ,.TP7D1 ( TP7D1 ) ,.TP7D0 ( TP7D0 )
 ,.TP6D3 ( TP6D3 ) ,.TP6D2 ( TP6D2 ) ,.TP6D1 ( TP6D1 ) ,.TP6D0 ( TP6D0 ) ,.TP5D3 ( TP5D3 ) ,.TP5D2 ( TP5D2 )
 ,.TP5D1 ( TP5D1 ) ,.TP5D0 ( TP5D0 ) ,.TP4D3 ( TP4D3 ) ,.TP4D2 ( TP4D2 ) ,.TP4D1 ( TP4D1 ) ,.TP4D0 ( TP4D0 )
 ,.TP3D3 ( TP3D3 ) ,.TP3D2 ( TP3D2 ) ,.TP3D1 ( TP3D1 ) ,.TP3D0 ( TP3D0 ) ,.TP2D3 ( TP2D3 ) ,.TP2D2 ( TP2D2 )
 ,.TP2D1 ( TP2D1 ) ,.TP2D0 ( TP2D0 ) ,.TP1D3 ( TP1D3 ) ,.TP1D2 ( TP1D2 ) ,.TP1D1 ( TP1D1 ) ,.TP1D0 ( TP1D0 )
 ,.TI11D3 ( TI11D3 ) ,.TI11D2 ( TI11D2 ) ,.TI11D1 ( TI11D1 ) ,.TI11D0 ( TI11D0 ) ,.TI10D3 ( TI10D3 ) ,.TI10D2 ( TI10D2 )
 ,.TI10D1 ( TI10D1 ) ,.TI10D0 ( TI10D0 ) ,.TI9D3 ( TI9D3 ) ,.TI9D2 ( TI9D2 ) ,.TI9D1 ( TI9D1 ) ,.TI9D0 ( TI9D0 )
 ,.TI8D3 ( TI8D3 ) ,.TI8D2 ( TI8D2 ) ,.TI8D1 ( TI8D1 ) ,.TI8D0 ( TI8D0 ) ,.TI7D3 ( TI7D3 ) ,.TI7D2 ( TI7D2 )
 ,.TI7D1 ( TI7D1 ) ,.TI7D0 ( TI7D0 ) ,.TI6D3 ( TI6D3 ) ,.TI6D2 ( TI6D2 ) ,.TI6D1 ( TI6D1 ) ,.TI6D0 ( TI6D0 )
 ,.TI5D3 ( TI5D3 ) ,.TI5D2 ( TI5D2 ) ,.TI5D1 ( TI5D1 ) ,.TI5D0 ( TI5D0 ) ,.TI4D3 ( TI4D3 ) ,.TI4D2 ( TI4D2 )
 ,.TI4D1 ( TI4D1 ) ,.TI4D0 ( TI4D0 ) ,.TI3D3 ( TI3D3 ) ,.TI3D2 ( TI3D2 ) ,.TI3D1 ( TI3D1 ) ,.TI3D0 ( TI3D0 )
 ,.TI2D3 ( TI2D3 ) ,.TI2D2 ( TI2D2 ) ,.TI2D1 ( TI2D1 ) ,.TI2D0 ( TI2D0 ) ,.TI1D3 ( TI1D3 ) ,.TI1D2 ( TI1D2 )
 ,.TI1D1 ( TI1D1 ) ,.TI1D0 ( TI1D0 ) ,.TI0D3 ( TI0D3 ) ,.TI0D2 ( TI0D2 ) ,.TI0D1 ( TI0D1 ) ,.TI0D0 ( TI0D0 )

  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/test.v
  TESTPIN ledtvdd_b (
   .ADDRH ( ADDRICE0 ) ,.EP ( ELEDTVDD_B ) ,.PIO ( UP ) ,.PUP ( DOWN ) ,.P ( LEDTVDD_B ) ,.TPD3 ( TI0D3 ) ,.TPD2 ( TI0D2 )
 ,.TPD1 ( TI0D1 ) ,.TPD0 ( TI0D0 ) ,.SYSRSOUTB ( SYSRSOUTB ) ,.ICEWR ( ICEWR ) ,.ICEDI0 ( ICEDI0 ) ,.ADDRPINRD ( ADDRPINRD )
 ,.ADDRPINMD ( ADDRPINMD ) ,.ADDRPINLV ( ADDRPINLV )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/test.v
  TESTPIN ledrun_b (
   .ADDRH ( ADDRICE1 ) ,.EP ( ELEDRUN_B ) ,.PIO ( UP ) ,.PUP ( DOWN ) ,.P ( LEDRUN_B ) ,.TPD3 ( TI1D3 ) ,.TPD2 ( TI1D2 )
 ,.TPD1 ( TI1D1 ) ,.TPD0 ( TI1D0 ) ,.SYSRSOUTB ( SYSRSOUTB ) ,.ICEWR ( ICEWR ) ,.ICEDI0 ( ICEDI0 ) ,.ADDRPINRD ( ADDRPINRD )
 ,.ADDRPINMD ( ADDRPINMD ) ,.ADDRPINLV ( ADDRPINLV )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/test.v
  TESTPIN ledreset_b (
   .ADDRH ( ADDRICE2 ) ,.EP ( ELEDRESET_B ) ,.PIO ( UP ) ,.PUP ( DOWN ) ,.P ( LEDRESET_B ) ,.TPD3 ( TI2D3 ) ,.TPD2 ( TI2D2 )
 ,.TPD1 ( TI2D1 ) ,.TPD0 ( TI2D0 ) ,.SYSRSOUTB ( SYSRSOUTB ) ,.ICEWR ( ICEWR ) ,.ICEDI0 ( ICEDI0 ) ,.ADDRPINRD ( ADDRPINRD )
 ,.ADDRPINMD ( ADDRPINMD ) ,.ADDRPINLV ( ADDRPINLV )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/test.v
  TESTPIN ledstandby_b (
   .ADDRH ( ADDRICE3 ) ,.EP ( ELEDSTANDBY_B ) ,.PIO ( UP ) ,.PUP ( DOWN ) ,.P ( LEDSTANDBY_B ) ,.TPD3 ( TI3D3 ) ,.TPD2 ( TI3D2 )
 ,.TPD1 ( TI3D1 ) ,.TPD0 ( TI3D0 ) ,.SYSRSOUTB ( SYSRSOUTB ) ,.ICEWR ( ICEWR ) ,.ICEDI0 ( ICEDI0 ) ,.ADDRPINRD ( ADDRPINRD )
 ,.ADDRPINMD ( ADDRPINMD ) ,.ADDRPINLV ( ADDRPINLV )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/test.v
  TESTPIN ledwait_b (
   .ADDRH ( ADDRICE4 ) ,.EP ( ELEDWAIT_B ) ,.PIO ( UP ) ,.PUP ( DOWN ) ,.P ( LEDWAIT_B ) ,.TPD3 ( TI4D3 ) ,.TPD2 ( TI4D2 )
 ,.TPD1 ( TI4D1 ) ,.TPD0 ( TI4D0 ) ,.SYSRSOUTB ( SYSRSOUTB ) ,.ICEWR ( ICEWR ) ,.ICEDI0 ( ICEDI0 ) ,.ADDRPINRD ( ADDRPINRD )
 ,.ADDRPINMD ( ADDRPINMD ) ,.ADDRPINLV ( ADDRPINLV )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/test.v
  TESTPIN ledclock_b (
   .ADDRH ( ADDRICE5 ) ,.EP ( ELEDCLOCK_B ) ,.PIO ( UP ) ,.PUP ( DOWN ) ,.P ( LEDCLOCK_B ) ,.TPD3 ( TI5D3 ) ,.TPD2 ( TI5D2 )
 ,.TPD1 ( TI5D1 ) ,.TPD0 ( TI5D0 ) ,.SYSRSOUTB ( SYSRSOUTB ) ,.ICEWR ( ICEWR ) ,.ICEDI0 ( ICEDI0 ) ,.ADDRPINRD ( ADDRPINRD )
 ,.ADDRPINMD ( ADDRPINMD ) ,.ADDRPINLV ( ADDRPINLV )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/test.v
  TESTPIN icesysres_b (
   .SYSRSOUTB ( ICESYSRES_B ) ,.ICEWR ( DOWN ) ,.ADDRH ( ADDRICE6 ) ,.EP ( EICESYSRES_B ) ,.PIO ( DOWN ) ,.PUP ( DOWN ) ,.P ( ICESYSRES_B )
 ,.TPD3 ( TI6D3 ) ,.TPD2 ( TI6D2 ) ,.TPD1 ( TI6D1 ) ,.TPD0 ( TI6D0 ) ,.ICEDI0 ( ICEDI0 ) ,.ADDRPINRD ( ADDRPINRD )
 ,.ADDRPINMD ( ADDRPINMD ) ,.ADDRPINLV ( ADDRPINLV )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/test.v
  TESTPIN icecpures_b (
   .ADDRH ( ADDRICE7 ) ,.EP ( EICECPURES_B ) ,.PIO ( DOWN ) ,.PUP ( DOWN ) ,.P ( ICECPURES_B ) ,.TPD3 ( TI7D3 ) ,.TPD2 ( TI7D2 )
 ,.TPD1 ( TI7D1 ) ,.TPD0 ( TI7D0 ) ,.SYSRSOUTB ( SYSRSOUTB ) ,.ICEWR ( ICEWR ) ,.ICEDI0 ( ICEDI0 ) ,.ADDRPINRD ( ADDRPINRD )
 ,.ADDRPINMD ( ADDRPINMD ) ,.ADDRPINLV ( ADDRPINLV )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/test.v
  TESTPIN eaconnect_b (
   .ADDRH ( ADDRICE8 ) ,.EP ( EEACONNECT_B ) ,.PIO ( DOWN ) ,.PUP ( DOWN ) ,.P ( EACONNECT_B ) ,.TPD3 ( TI8D3 ) ,.TPD2 ( TI8D2 )
 ,.TPD1 ( TI8D1 ) ,.TPD0 ( TI8D0 ) ,.SYSRSOUTB ( SYSRSOUTB ) ,.ICEWR ( ICEWR ) ,.ICEDI0 ( ICEDI0 ) ,.ADDRPINRD ( ADDRPINRD )
 ,.ADDRPINMD ( ADDRPINMD ) ,.ADDRPINLV ( ADDRPINLV )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/test.v
  TESTPIN tcconnect_b (
   .ADDRH ( ADDRICE9 ) ,.EP ( ETCCONNECT_B ) ,.PIO ( DOWN ) ,.PUP ( DOWN ) ,.P ( TCCONNECT_B ) ,.TPD3 ( TI9D3 ) ,.TPD2 ( TI9D2 )
 ,.TPD1 ( TI9D1 ) ,.TPD0 ( TI9D0 ) ,.SYSRSOUTB ( SYSRSOUTB ) ,.ICEWR ( ICEWR ) ,.ICEDI0 ( ICEDI0 ) ,.ADDRPINRD ( ADDRPINRD )
 ,.ADDRPINMD ( ADDRPINMD ) ,.ADDRPINLV ( ADDRPINLV )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/test.v
  TESTPIN tvddon (
   .ADDRH ( ADDRICE10 ) ,.EP ( ETVDDON ) ,.PIO ( DOWN ) ,.PUP ( DOWN ) ,.P ( TVDDON ) ,.TPD3 ( TI10D3 ) ,.TPD2 ( TI10D2 )
 ,.TPD1 ( TI10D1 ) ,.TPD0 ( TI10D0 ) ,.SYSRSOUTB ( SYSRSOUTB ) ,.ICEWR ( ICEWR ) ,.ICEDI0 ( ICEDI0 ) ,.ADDRPINRD ( ADDRPINRD )
 ,.ADDRPINMD ( ADDRPINMD ) ,.ADDRPINLV ( ADDRPINLV )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/test.v
  TESTPIN tvddsel (
   .ADDRH ( ADDRICE11 ) ,.EP ( ETVDDSEL ) ,.PIO ( UP ) ,.PUP ( DOWN ) ,.P ( TVDDSELB ) ,.TPD3 ( TI11D3 ) ,.TPD2 ( TI11D2 )
 ,.TPD1 ( TI11D1 ) ,.TPD0 ( TI11D0 ) ,.SYSRSOUTB ( SYSRSOUTB ) ,.ICEWR ( ICEWR ) ,.ICEDI0 ( ICEDI0 ) ,.ADDRPINRD ( ADDRPINRD )
 ,.ADDRPINMD ( ADDRPINMD ) ,.ADDRPINLV ( ADDRPINLV )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/ice_other.v
  ice_other ice_other (
   .UP ( UP ) ,.DOWN ( DOWN ) ,.TVDDSELB ( TVDDSELB ) ,.TVDDSEL ( TVDDSEL ) ,.EROMWAIT ( EROMWAIT ) ,.TMEMWAIT ( TMEMWAIT ) ,.WAITOR ( WAITOR )
 ,.CLK30MHZ ( CLK30MHZ ) ,.CLK30MHZ_GB ( CLK30MHZ_GB ) ,.ICEDI_PRE31 ( ICEDI_PRE31 ) ,.ICEDI_PRE23 ( ICEDI_PRE23 ) ,.ICEDI_PRE15 ( ICEDI_PRE15 ) ,.ICEDI_PRE30 ( ICEDI_PRE30 )
 ,.ICEDI_PRE22 ( ICEDI_PRE22 ) ,.ICEDI_PRE14 ( ICEDI_PRE14 ) ,.ICEDI_PRE29 ( ICEDI_PRE29 ) ,.ICEDI_PRE28 ( ICEDI_PRE28 ) ,.ICEDI_PRE27 ( ICEDI_PRE27 ) ,.ICEDI_PRE19 ( ICEDI_PRE19 )
 ,.ICEDI_PRE26 ( ICEDI_PRE26 ) ,.ICEDI_PRE18 ( ICEDI_PRE18 ) ,.ICEDI_PRE25 ( ICEDI_PRE25 ) ,.ICEDI_PRE17 ( ICEDI_PRE17 ) ,.ICEDI_PRE24 ( ICEDI_PRE24 ) ,.ICEDI_PRE16 ( ICEDI_PRE16 )
 ,.ICEDI_PRE21 ( ICEDI_PRE21 ) ,.ICEDI_PRE13 ( ICEDI_PRE13 ) ,.ICEDI_PRE20 ( ICEDI_PRE20 ) ,.ICEDI_PRE12 ( ICEDI_PRE12 ) ,.ICEDI_PRE11 ( ICEDI_PRE11 ) ,.ICEDI_PRE10 ( ICEDI_PRE10 )
 ,.ICEDI_PRE9 ( ICEDI_PRE9 ) ,.ICEDI_PRE8 ( ICEDI_PRE8 ) ,.ICEDI_PRE7 ( ICEDI_PRE7 ) ,.ICEDI_PRE6 ( ICEDI_PRE6 ) ,.ICEDI_PRE5 ( ICEDI_PRE5 ) ,.ICEDI_PRE4 ( ICEDI_PRE4 )
 ,.ICEDI_PRE3 ( ICEDI_PRE3 ) ,.ICEDI_PRE2 ( ICEDI_PRE2 ) ,.ICEDI_PRE1 ( ICEDI_PRE1 ) ,.ETVDDSEL ( ETVDDSEL ) ,.ELEDTVDD_B ( ELEDTVDD_B ) ,.ELEDCLOCK_B ( ELEDCLOCK_B )
 ,.ELEDRUN_B ( ELEDRUN_B ) ,.ELEDRESET_B ( ELEDRESET_B ) ,.ELEDSTANDBY_B ( ELEDSTANDBY_B ) ,.ELEDWAIT_B ( ELEDWAIT_B ) ,.ICECPURES_B ( ICECPURES_B ) ,.TCCONNECT_B ( TCCONNECT_B )
 ,.EACONNECT_B ( EACONNECT_B ) ,.TVDDON ( TVDDON ) ,.ICERD_PRE ( ICERD_PRE ) ,.EXMAPOUT ( EXMAPOUT ) ,.ICEIFA_PRE1 ( ICEIFA_PRE1 ) ,.ICEIFA_PRE0 ( ICEIFA_PRE0 )
 ,.ICEFLERRC ( ICEFLERRC ) ,.ICEFLERRD ( ICEFLERRD ) ,.ICEFLERR ( ICEFLERR )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacroSuite/ICEMacro/trunk/Source/DFlashEmu1.v
  DFLASHEMU1 dflashemu (
   .CLK30MHZ ( CLK30MHZ_GB ) ,.CLK60MHZ ( CLK60MHZ ) ,.DRDCLKP1_OUT ( DRDCLKP1_OUT ) ,.DWWR_OUT ( DWWR_OUT ) ,.DCER_OUT ( DCER_OUT ) ,.DSER_OUT ( DSER_OUT ) ,.DMRG00_OUT ( DMRG00_OUT )
 ,.DMRG01_OUT ( DMRG01_OUT ) ,.DMRG10_OUT ( DMRG10_OUT ) ,.DMRG11_OUT ( DMRG11_OUT ) ,.DMRG12_OUT ( DMRG12_OUT ) ,.DDIS_OUT ( DDIS_OUT ) ,.ICEDOU30 ( ICEDOU30 )
 ,.ICEDOU22 ( ICEDOU22 ) ,.ICEDOU14 ( ICEDOU14 ) ,.DREAD_OUT ( DREAD_OUT ) ,.DFCLK_OUT ( DFCLK_OUT ) ,.ICEIFA31 ( ICEIFA31 ) ,.ICEIFA23 ( ICEIFA23 )
 ,.ICEIFA15 ( ICEIFA15 ) ,.ICEIFA30 ( ICEIFA30 ) ,.ICEIFA22 ( ICEIFA22 ) ,.ICEIFA14 ( ICEIFA14 ) ,.ICEIFA29 ( ICEIFA29 ) ,.ICEIFA28 ( ICEIFA28 )
 ,.ICEIFA27 ( ICEIFA27 ) ,.ICEIFA19 ( ICEIFA19 ) ,.ICEIFA26 ( ICEIFA26 ) ,.ICEIFA18 ( ICEIFA18 ) ,.ICEIFA25 ( ICEIFA25 ) ,.ICEIFA17 ( ICEIFA17 )
 ,.ICEIFA24 ( ICEIFA24 ) ,.ICEIFA16 ( ICEIFA16 ) ,.ICEIFA21 ( ICEIFA21 ) ,.ICEIFA13 ( ICEIFA13 ) ,.ICEIFA20 ( ICEIFA20 ) ,.ICEIFA12 ( ICEIFA12 )
 ,.ICEIFA11 ( ICEIFA11 ) ,.ICEIFA10 ( ICEIFA10 ) ,.ICEIFA9 ( ICEIFA9 ) ,.ICEIFA8 ( ICEIFA8 ) ,.ICEIFA7 ( ICEIFA7 ) ,.ICEIFA6 ( ICEIFA6 )
 ,.ICEIFA5 ( ICEIFA5 ) ,.ICEIFA4 ( ICEIFA4 ) ,.ICEIFA3 ( ICEIFA3 ) ,.ICEIFA2 ( ICEIFA2 ) ,.ICEIFA1 ( ICEIFA1 ) ,.ICEIFA0 ( ICEIFA0 )
 ,.ICEDOU31 ( ICEDOU31 ) ,.ICEDOU23 ( ICEDOU23 ) ,.ICEDOU15 ( ICEDOU15 ) ,.ICEDOU29 ( ICEDOU29 ) ,.ICEDOU28 ( ICEDOU28 ) ,.ICEDOU27 ( ICEDOU27 )
 ,.ICEDOU19 ( ICEDOU19 ) ,.ICEDOU26 ( ICEDOU26 ) ,.ICEDOU18 ( ICEDOU18 ) ,.ICEDOU25 ( ICEDOU25 ) ,.ICEDOU17 ( ICEDOU17 ) ,.ICEDOU24 ( ICEDOU24 )
 ,.ICEDOU16 ( ICEDOU16 ) ,.ICEDOU21 ( ICEDOU21 ) ,.ICEDOU13 ( ICEDOU13 ) ,.ICEDOU20 ( ICEDOU20 ) ,.ICEDOU12 ( ICEDOU12 ) ,.ICEDOU11 ( ICEDOU11 )
 ,.ICEDOU10 ( ICEDOU10 ) ,.ICEDOU9 ( ICEDOU9 ) ,.ICEDOU8 ( ICEDOU8 ) ,.ICEDOU7 ( ICEDOU7 ) ,.ICEDOU6 ( ICEDOU6 ) ,.ICEDOU5 ( ICEDOU5 )
 ,.ICEDOU4 ( ICEDOU4 ) ,.ICEDOU3 ( ICEDOU3 ) ,.ICEDOU2 ( ICEDOU2 ) ,.ICEDOU1 ( ICEDOU1 ) ,.ICEDOU0 ( ICEDOU0 ) ,.ICEDI31 ( ICEDI31 )
 ,.ICEDI23 ( ICEDI23 ) ,.ICEDI15 ( ICEDI15 ) ,.ICEDI30 ( ICEDI30 ) ,.ICEDI22 ( ICEDI22 ) ,.ICEDI14 ( ICEDI14 ) ,.ICEDI29 ( ICEDI29 )
 ,.ICEDI28 ( ICEDI28 ) ,.ICEDI27 ( ICEDI27 ) ,.ICEDI19 ( ICEDI19 ) ,.ICEDI26 ( ICEDI26 ) ,.ICEDI18 ( ICEDI18 ) ,.ICEDI25 ( ICEDI25 )
 ,.ICEDI17 ( ICEDI17 ) ,.ICEDI24 ( ICEDI24 ) ,.ICEDI16 ( ICEDI16 ) ,.ICEDI21 ( ICEDI21 ) ,.ICEDI13 ( ICEDI13 ) ,.ICEDI20 ( ICEDI20 )
 ,.ICEDI12 ( ICEDI12 ) ,.ICEDI11 ( ICEDI11 ) ,.ICEDI10 ( ICEDI10 ) ,.ICEDI9 ( ICEDI9 ) ,.ICEDI8 ( ICEDI8 ) ,.ICEDI7 ( ICEDI7 )
 ,.ICEDI6 ( ICEDI6 ) ,.ICEDI5 ( ICEDI5 ) ,.ICEDI4 ( ICEDI4 ) ,.ICEDI3 ( ICEDI3 ) ,.ICEDI2 ( ICEDI2 ) ,.ICEDI1 ( ICEDI1 )
 ,.ICEDI0 ( ICEDI0 ) ,.ICEWR ( ICEWR ) ,.SVMOD ( SVMOD ) ,.SVMODF ( SVMODF ) ,.ALT1 ( ALT1 ) ,.PREFIX ( PREFIX )
 ,.SLFLASH ( SLFLASH ) ,.FLREAD ( FLREAD ) ,.PA19 ( PA19 ) ,.FCLK ( FCLK ) ,.PA18 ( PA18 ) ,.PA17 ( PA17 )
 ,.PA16 ( PA16 ) ,.PA15 ( PA15 ) ,.PA14 ( PA14 ) ,.PA13 ( PA13 ) ,.PA12 ( PA12 ) ,.PA11 ( PA11 )
 ,.PA10 ( PA10 ) ,.PA9 ( PA9 ) ,.PA8 ( PA8 ) ,.PA7 ( PA7 ) ,.PA6 ( PA6 ) ,.PA5 ( PA5 )
 ,.DW9 ( DW9 ) ,.PA4 ( PA4 ) ,.DW8 ( DW8 ) ,.PA3 ( PA3 ) ,.DW7 ( DW7 ) ,.PA2 ( PA2 )
 ,.DW6 ( DW6 ) ,.SLMEM ( SLMEM ) ,.EXMA3 ( EXMA3 ) ,.EXMA2 ( EXMA2 ) ,.EXMA1 ( EXMA1 ) ,.EXMA0 ( EXMA0 )
 ,.MA15 ( MA15 ) ,.MA14 ( MA14 ) ,.MA13 ( MA13 ) ,.MA12 ( MA12 ) ,.BEU2 ( BEU2 ) ,.MA11 ( MA11 )
 ,.BEU1 ( BEU1 ) ,.MA10 ( MA10 ) ,.BEU0 ( BEU0 ) ,.MA9 ( MA9 ) ,.DW1 ( DW1 ) ,.MA8 ( MA8 )
 ,.DW0 ( DW0 ) ,.MA7 ( MA7 ) ,.MA6 ( MA6 ) ,.MA5 ( MA5 ) ,.MA4 ( MA4 ) ,.MA3 ( MA3 )
 ,.MA2 ( MA2 ) ,.MA1 ( MA1 ) ,.MA0 ( MA0 ) ,.MDW15 ( MDW15 ) ,.MDW14 ( MDW14 ) ,.MDW13 ( MDW13 )
 ,.MDW12 ( MDW12 ) ,.MDW11 ( MDW11 ) ,.MDW10 ( MDW10 ) ,.MDW9 ( MDW9 ) ,.MDW8 ( MDW8 ) ,.MDW7 ( MDW7 )
 ,.MDW6 ( MDW6 ) ,.MDW5 ( MDW5 ) ,.MDW4 ( MDW4 ) ,.MDW3 ( MDW3 ) ,.MDW2 ( MDW2 ) ,.MDW1 ( MDW1 )
 ,.MDW0 ( MDW0 ) ,.DFMDR15 ( DFMDR15 ) ,.DFMDR14 ( DFMDR14 ) ,.DFMDR13 ( DFMDR13 ) ,.DFMDR12 ( DFMDR12 ) ,.DFMDR11 ( DFMDR11 )
 ,.DFMDR10 ( DFMDR10 ) ,.DFMDR9 ( DFMDR9 ) ,.DFMDR8 ( DFMDR8 ) ,.DFMDR7 ( DFMDR7 ) ,.DFMDR6 ( DFMDR6 ) ,.DFMDR5 ( DFMDR5 )
 ,.DFMDR4 ( DFMDR4 ) ,.DFMDR3 ( DFMDR3 ) ,.DFMDR2 ( DFMDR2 ) ,.DFMDR1 ( DFMDR1 ) ,.DFMDR0 ( DFMDR0 ) ,.CPUWR ( CPUWR )
 ,.CPURD ( CPURD ) ,.WDOP ( WDOP ) ,.SLBMEM ( SLBMEM ) ,.DCLKSEL1 ( DCLKSEL1 ) ,.DRDCLK ( DRDCLK ) ,.DRDCLKC1 ( DRDCLKC1 )
 ,.RDCLKP1 ( RDCLKP1 ) ,.DCE0 ( DCE0 ) ,.AF19 ( AF19 ) ,.AF18 ( AF18 ) ,.AF17 ( AF17 ) ,.DA13 ( DA13 )
 ,.AF16 ( AF16 ) ,.DA12 ( DA12 ) ,.AF15 ( AF15 ) ,.DA11 ( DA11 ) ,.AF14 ( AF14 ) ,.DA10 ( DA10 )
 ,.AF13 ( AF13 ) ,.AF12 ( AF12 ) ,.AF11 ( AF11 ) ,.AF10 ( AF10 ) ,.AF9 ( AF9 ) ,.DA7 ( DA7 )
 ,.AF8 ( AF8 ) ,.DA6 ( DA6 ) ,.AF7 ( AF7 ) ,.DA5 ( DA5 ) ,.AF6 ( AF6 ) ,.DA4 ( DA4 )
 ,.AF5 ( AF5 ) ,.DA3 ( DA3 ) ,.AF4 ( AF4 ) ,.DA2 ( DA2 ) ,.AF3 ( AF3 ) ,.DA1 ( DA1 )
 ,.AF2 ( AF2 ) ,.DA0 ( DA0 ) ,.AF1 ( AF1 ) ,.AF0 ( AF0 ) ,.DA9 ( DA9 ) ,.DA8 ( DA8 )
 ,.DRO11 ( DRO11 ) ,.DRO10 ( DRO10 ) ,.DRO9 ( DRO9 ) ,.DRO8 ( DRO8 ) ,.DRO7 ( DRO7 ) ,.DRO6 ( DRO6 )
 ,.DRO5 ( DRO5 ) ,.DRO4 ( DRO4 ) ,.DRO3 ( DRO3 ) ,.DRO2 ( DRO2 ) ,.DRO1 ( DRO1 ) ,.DRO0 ( DRO0 )
 ,.DWWR ( DWWR ) ,.DCER ( DCER ) ,.DSER ( DSER ) ,.DMRG00 ( DMRG00 ) ,.DMRG01 ( DMRG01 ) ,.DMRG10 ( DMRG10 )
 ,.DMRG11 ( DMRG11 ) ,.DMRG12 ( DMRG12 ) ,.DDIS ( DDIS ) ,.DREAD ( DREAD ) ,.DWED ( DWED ) ,.PROGI ( PROGI )
 ,.DW11 ( DW11 ) ,.DW10 ( DW10 ) ,.DW5 ( DW5 ) ,.DW4 ( DW4 ) ,.DW3 ( DW3 ) ,.DW2 ( DW2 )
 ,.ICEFLERRD ( ICEFLERRD ) ,.CPURSOUTB ( CPURSOUTB ) ,.SYSRSOUTB ( SYSRSOUTB ) ,.BASECK ( BASECK )
  ) ;
endmodule


// $Id: idversion.v,v 1.6 2007-10-03 04:02:52 tsuno3 Exp $
// v1.7 : Add FNAVAIL emulation register.
//        And TIMER block 32MHz available.

module IDVERSION (
	IDVER31, IDVER30, IDVER29, IDVER28,
	IDVER27, IDVER26, IDVER25, IDVER24,
	IDVER23, IDVER22, IDVER21, IDVER20,
	IDVER19, IDVER18, IDVER17, IDVER16,
	IDVER15, IDVER14, IDVER13, IDVER12,
	IDVER11, IDVER10, IDVER9, IDVER8,
	IDVER7, IDVER6, IDVER5, IDVER4,
	IDVER3, IDVER2, IDVER1, IDVER0,
	ICEIFA31, ICEIFA30, ICEIFA29, ICEIFA28,
	ICEIFA27, ICEIFA26, ICEIFA25, ICEIFA24,
	ICEIFA23, ICEIFA22, ICEIFA21, ICEIFA20,
	ICEIFA19, ICEIFA18, ICEIFA17, ICEIFA16,
	ICEIFA15, ICEIFA14, ICEIFA13, ICEIFA12,
	ICEIFA11, ICEIFA10, ICEIFA9, ICEIFA8,
	ICEIFA7, ICEIFA6, ICEIFA5, ICEIFA4,
	ICEIFA3, ICEIFA2, ICEIFA1, ICEIFA0,
	ICEDO31, ICEDO30, ICEDO29, ICEDO28,
	ICEDO27, ICEDO26, ICEDO25, ICEDO24,
	ICEDO23, ICEDO22, ICEDO21, ICEDO20,
	ICEDO19, ICEDO18, ICEDO17, ICEDO16,
	ICEDO15, ICEDO14, ICEDO13, ICEDO12,
	ICEDO11, ICEDO10, ICEDO9, ICEDO8,
	ICEDO7, ICEDO6, ICEDO5, ICEDO4,
	ICEDO3, ICEDO2, ICEDO1, ICEDO0
);
	input	IDVER31, IDVER30, IDVER29, IDVER28,
			IDVER27, IDVER26, IDVER25, IDVER24,
			IDVER23, IDVER22, IDVER21, IDVER20,
			IDVER19, IDVER18, IDVER17, IDVER16,
			IDVER15, IDVER14, IDVER13, IDVER12,
			IDVER11, IDVER10, IDVER9, IDVER8,
			IDVER7, IDVER6, IDVER5, IDVER4,
			IDVER3, IDVER2, IDVER1, IDVER0;
	input	ICEIFA31, ICEIFA30, ICEIFA29, ICEIFA28,
			ICEIFA27, ICEIFA26, ICEIFA25, ICEIFA24,
			ICEIFA23, ICEIFA22, ICEIFA21, ICEIFA20,
			ICEIFA19, ICEIFA18, ICEIFA17, ICEIFA16,
			ICEIFA15, ICEIFA14, ICEIFA13, ICEIFA12,
			ICEIFA11, ICEIFA10, ICEIFA9, ICEIFA8,
			ICEIFA7, ICEIFA6, ICEIFA5, ICEIFA4,
			ICEIFA3, ICEIFA2, ICEIFA1, ICEIFA0;
	output	ICEDO31, ICEDO30, ICEDO29, ICEDO28,
			ICEDO27, ICEDO26, ICEDO25, ICEDO24,
			ICEDO23, ICEDO22, ICEDO21, ICEDO20,
			ICEDO19, ICEDO18, ICEDO17, ICEDO16,
			ICEDO15, ICEDO14, ICEDO13, ICEDO12,
			ICEDO11, ICEDO10, ICEDO9, ICEDO8,
			ICEDO7, ICEDO6, ICEDO5, ICEDO4,
			ICEDO3, ICEDO2, ICEDO1, ICEDO0;
	
	wire [31:0] IDVER, ICEDO;
	wire sel_idver;

	assign	{
		ICEDO31, ICEDO30, ICEDO29, ICEDO28, ICEDO27, ICEDO26, ICEDO25, ICEDO24,
		ICEDO23, ICEDO22, ICEDO21, ICEDO20, ICEDO19, ICEDO18, ICEDO17, ICEDO16,
		ICEDO15, ICEDO14, ICEDO13, ICEDO12, ICEDO11, ICEDO10, ICEDO9, ICEDO8,
		ICEDO7, ICEDO6, ICEDO5, ICEDO4, ICEDO3, ICEDO2, ICEDO1, ICEDO0
	} = ICEDO;
	assign	IDVER = {
		IDVER31, IDVER30, IDVER29, IDVER28, IDVER27, IDVER26, IDVER25, IDVER24,
		IDVER23, IDVER22, IDVER21, IDVER20, IDVER19, IDVER18, IDVER17, IDVER16,
		IDVER15, IDVER14, IDVER13, IDVER12, IDVER11, IDVER10, IDVER9, IDVER8,
		IDVER7, IDVER6, IDVER5, IDVER4, IDVER3, IDVER2, IDVER1, IDVER0
	};
	wire [31:0] iceifa = {
		ICEIFA31, ICEIFA30, ICEIFA29, ICEIFA28, ICEIFA27, ICEIFA26, ICEIFA25, ICEIFA24,
		ICEIFA23, ICEIFA22, ICEIFA21, ICEIFA20, ICEIFA19, ICEIFA18, ICEIFA17, ICEIFA16,
		ICEIFA15, ICEIFA14, ICEIFA13, ICEIFA12, ICEIFA11, ICEIFA10, ICEIFA9, ICEIFA8,
		ICEIFA7,  ICEIFA6,  ICEIFA5,  ICEIFA4,  ICEIFA3,  ICEIFA2,  ICEIFA1, ICEIFA0
	};
	assign sel_idver   = iceifa[27] & iceifa[23] & iceifa[15] ;                               // 0880_8xxxH : IDVER
	assign sel_fnavail = iceifa[27] & iceifa[23] & iceifa[14] & { iceifa[11:0] == 12'h008 } ; // 0880_4008H : FNAVAIL

	assign ICEDO = (sel_idver)   ? IDVER :
                       (sel_fnavail) ? {32'b0000_0000_0000_0000__0000_0000_0000_0011} :
  		                        // bit31-2 : Unused
		                        // bit1 : TIMER block 32MHz available
		                        // bit0 : TIMETAG block 32MHz available
                       32'h0000_0000 ;

endmodule

//  file name   ... /proj/78k0r_11/78k0r_kx4/_ice/_make_chip/_eva_top/_library/eva_top_056.v
//  top module  ... /proj/78k0r_11/78k0r_kx4/_ice/_make_chip/_eva_top/_library/eva_top_056.v EVA_TOP
//  version     ... 1.00
//  designer    ... T.Tsunoda
//  refer to    ... make_chip.para
 
module EVA_TOP (
  CLK30MHZ ,EVAOSCMCLK ,RESET_B ,ICESYSRES_B ,ICECPURES_B ,EACONNECT_B ,TCCONNECT_B ,TVDDSEL ,TVDDON ,LEDCLOCK_B ,LEDRESET_B 
 ,LEDRUN_B ,LEDSTANDBY_B ,LEDTVDD_B ,LEDWAIT_B ,USBCLK ,USBRD_B ,USBWR0_B ,USBWAIT_B ,USBA1 ,USBA2
 ,PPUP0 ,USBA3 ,PPUP1 ,USBA4 ,PPUP2 ,USBA19 ,PPUP15 ,PPUP31 ,USBA20 ,USBA21
 ,USBD0 ,PPUP4 ,USBD1 ,PPUP5 ,USBD2 ,PPUP6 ,USBD3 ,PPUP7 ,USBD4 ,PPUP8
 ,USBD5 ,PPUP9 ,USBD6 ,USBD7 ,USBD8 ,USBD9 ,USBD10 ,PPUP18 ,PPUP26 ,USBD11
 ,PPUP19 ,PPUP27 ,USBD12 ,PPUP28 ,USBD13 ,PPUP29 ,USBD14 ,USBD15 ,EROMCLK ,EROMCSB
 ,EROMPA2 ,EROMWRB ,EROMRDB ,EROMPA0 ,EROMPA1 ,EROMPA3 ,EROMPA4 ,EROMPA5 ,EROMPA6 ,EROMPD0
 ,EROMPA7 ,EROMPD1 ,EROMPA8 ,EROMPD2 ,EROMPA9 ,EROMPD3 ,EROMPA10 ,EROMPA11 ,EROMPA12 ,EROMPA13
 ,EROMPA14 ,EROMPA15 ,EROMPA16 ,EROMPA17 ,EROMPD4 ,EROMPD5 ,EROMPD6 ,EROMPD7 ,EROMPD8 ,EROMPD9
 ,EROMPD10 ,EROMPD11 ,EROMPD12 ,EROMPD20 ,EROMPD13 ,EROMPD21 ,EROMPD14 ,EROMPD22 ,EROMPD30 ,EROMPD15
 ,EROMPD23 ,EROMPD31 ,EROMPD16 ,EROMPD24 ,EROMPD32 ,EROMPD17 ,EROMPD25 ,EROMPD33 ,EROMPD18 ,EROMPD26
 ,EROMPD34 ,EROMPD19 ,EROMPD27 ,EROMPD35 ,EROMPD28 ,EROMPD29 ,DIS_OUT ,WWR_OUT ,MRG00_OUT ,MRG01_OUT
 ,MRG10_OUT ,MRG11_OUT ,MRG12_OUT ,READ_OUT ,FCLK_OUT ,RDCLKP1_OUT ,PROGI_OUT ,CER_OUT ,SER_OUT ,EXA_OUT
 ,EXER_OUT ,BFA_OUT ,TMEMCLK0 ,TMEMCLK1 ,TMEMCLK2 ,TMEMCS_B ,TMEMRD_B ,TMEMWR_B ,TMEMA0 ,TMEMA1
 ,TMEMA2 ,TMEMA3 ,TMEMA4 ,TMEMA5 ,TMEMA6 ,TMEMD0 ,TMEMA7 ,TMEMD1 ,TMEMA8 ,TMEMD2
 ,TMEMA9 ,TMEMD3 ,TMEMA10 ,TMEMA11 ,TMEMA12 ,TMEMA13 ,TMEMA14 ,TMEMA15 ,TMEMA16 ,TMEMD4
 ,TMEMD5 ,TMEMD6 ,TMEMD7 ,TMEMD8 ,TMEMD9 ,TMEMD10 ,TMEMD11 ,TMEMD12 ,TMEMD20 ,TMEMD13
 ,TMEMD21 ,TMEMD14 ,TMEMD22 ,TMEMD30 ,TMEMD15 ,TMEMD23 ,TMEMD31 ,TMEMD16 ,TMEMD24 ,TMEMD32
 ,TMEMD40 ,TMEMD17 ,TMEMD25 ,TMEMD33 ,TMEMD41 ,TMEMD18 ,TMEMD26 ,TMEMD34 ,TMEMD42 ,TMEMD50
 ,TMEMD19 ,TMEMD27 ,TMEMD35 ,TMEMD43 ,TMEMD51 ,TMEMD28 ,TMEMD36 ,TMEMD44 ,TMEMD52 ,TMEMD60
 ,TMEMD29 ,TMEMD37 ,TMEMD45 ,TMEMD53 ,TMEMD61 ,TMEMD38 ,TMEMD46 ,TMEMD54 ,TMEMD62 ,TMEMD70
 ,TMEMD39 ,TMEMD47 ,TMEMD55 ,TMEMD63 ,TMEMD71 ,TMEMD48 ,TMEMD56 ,TMEMD64 ,TMEMD72 ,TMEMD80
 ,TMEMD49 ,TMEMD57 ,TMEMD65 ,TMEMD73 ,TMEMD81 ,TMEMD58 ,TMEMD66 ,TMEMD74 ,TMEMD82 ,TMEMD90
 ,TMEMD59 ,TMEMD67 ,TMEMD75 ,TMEMD83 ,TMEMD91 ,TMEMD68 ,TMEMD76 ,TMEMD84 ,TMEMD92 ,TMEMD69
 ,TMEMD77 ,TMEMD85 ,TMEMD93 ,TMEMD78 ,TMEMD86 ,TMEMD94 ,TMEMD79 ,TMEMD87 ,TMEMD95 ,TMEMD88
 ,TMEMD96 ,TMEMD89 ,TMEMD97 ,TMEMD98 ,TMEMD99 ,TMEMD100 ,TMEMD101 ,TMEMD102 ,TMEMD103 ,TMEMD104
 ,TMEMD105 ,TMEMD106 ,TMEMD107 ,LVISEL ,P121 ,P122 ,P130 ,AP10 ,P123 ,AP11
 ,P124 ,P140 ,AP12 ,AP20 ,P00 ,P01 ,P02 ,P10 ,P03 ,P11
 ,PTTL03 ,PTTL11 ,P04 ,P12 ,P20 ,PTTL04 ,P05 ,P13 ,P21 ,AP1
 ,P06 ,P14 ,P22 ,P30 ,AP2 ,PTTL10 ,PTTL13 ,PTTL14 ,P15 ,P23
 ,P31 ,AP3 ,PTTL15 ,P16 ,P24 ,P40 ,AP4 ,PTTL16 ,P17 ,P25
 ,P41 ,AP5 ,PTTL17 ,P26 ,P42 ,P50 ,AP6 ,P27 ,P43 ,P51
 ,AP7 ,P52 ,P60 ,AP8 ,P53 ,P61 ,AP9 ,P54 ,P62 ,P70
 ,P55 ,P63 ,P71 ,P72 ,P73 ,P74 ,P75 ,P76 ,P77 ,P120
 ,P137 ,AP17 ,AP25 ,AP33 ,AP41 ,P141 ,AP13 ,AP21 ,P146 ,AP18
 ,AP26 ,AP34 ,AP42 ,AP50 ,P147 ,AP19 ,AP27 ,AP35 ,AP43 ,AP51
 ,PPUP3 ,PPUP10 ,PPUP11 ,PPUP12 ,PPUP20 ,PPUP13 ,PPUP21 ,PPUP14 ,PPUP30 ,PPUP16
 ,PPUP24 ,PPUP17 ,PPUP25 ,PUPLE0 ,PUPLE1 ,PUPLE2 ,PUPLE3 ,PUPLE4 ,PUPLE5 ,PSSC0
 ,PSSC1 ,PSSC2 ,PSSC3 ,PSSC4 ,PSSC5 ,PIO00 ,PIO01 ,PIO02 ,PIO10 ,PIO03
 ,PIO11 ,PIO04 ,PIO12 ,PIO20 ,PIO05 ,PIO13 ,PIO21 ,PIO06 ,PIO14 ,PIO22
 ,PIO30 ,PIO15 ,PIO23 ,PIO31 ,PIO16 ,PIO24 ,PIO40 ,PIO17 ,PIO25 ,PIO41
 ,PIO26 ,PIO42 ,PIO50 ,PIO27 ,PIO43 ,PIO51 ,PIO52 ,PIO60 ,PIO53 ,PIO61
 ,PIO54 ,PIO62 ,PIO70 ,PIO55 ,PIO63 ,PIO71 ,PIO72 ,PIO73 ,PIO74 ,PIO75
 ,PIO76 ,PIO77 ,PIO120 ,PIO121 ,PIO122 ,PIO130 ,PIO123 ,PIO124 ,PIO140 ,PIO141
 ,PIO146 ,PIO147 ,ADINT_B ,AD_DB9 ,AD_DB8 ,AD_DB7 ,AD_DB6 ,AD_DB5 ,AD_DB4 ,AD_DB3
 ,AD_DB2 ,AD_DB1 ,AD_DB0 ,ADCS_B ,ADRD_B ,ADSH_B ,AD_A4 ,AD_A3 ,AD_A2 ,AD_A1
 ,AD_A0 ,ADGSELMOD ,PORTEN_B0 ,PORTEN_B1 ,PORTEN_B2 ,PORTEN_B3 ,PORTEN_B4 ,PORTEN_B5 ,PORTEN_B6 ,PORTEN_B7
 ,PORTEN_B8 ,PORTEN_B9 ,PORTEN_B10 ,PORTEN_B11 ,EMVDDSEL_B ,ADVSELMOD ,AP14 ,AP22 ,AP30 ,AP15
 ,AP23 ,AP31 ,AP16 ,AP24 ,AP32 ,AP40 ,AP28 ,AP36 ,AP44 ,AP52
 ,AP60 ,AP29 ,AP37 ,AP45 ,AP53 ,AP61 ,AP38 ,AP46 ,AP54 ,AP62
 ,AP39 ,AP47 ,AP55 ,AP63 ,AP48 ,AP56 ,AP64 ,AP49 ,AP57 ,AP65
 ,AP58 ,AP59 ,APIO1 ,APIO2 ,APIO3 ,APIO4 ,APIO5 ,APIO6 ,APIO7 ,APIO8
 ,APIO9 ,APIO10 ,APIO11 ,APIO12 ,APIO20 ,APIO13 ,APIO21 ,APIO14 ,APIO22 ,APIO30
 ,APIO15 ,APIO23 ,APIO31 ,APIO16 ,APIO24 ,APIO32 ,APIO40 ,APIO17 ,APIO25 ,APIO33
 ,APIO41 ,APIO18 ,APIO26 ,APIO34 ,APIO42 ,APIO50 ,APIO19 ,APIO27 ,APIO35 ,APIO43
 ,APIO51 ,APIO28 ,APIO36 ,APIO44 ,APIO52 ,APIO60 ,APIO29 ,APIO37 ,APIO45 ,APIO53
 ,APIO61 ,APIO38 ,APIO46 ,APIO54 ,APIO62 ,APIO39 ,APIO47 ,APIO55 ,APIO63 ,APIO48
 ,APIO56 ,APIO64 ,APIO49 ,APIO57 ,APIO65 ,APIO58 ,APIO59 ,PIO_ANALOG0 ,PIO_ANALOG1 ,PIO_ANALOG2
 ,PIO_ANALOG3 ,PIO_ANALOG4 ,PIO_ANALOG5 ,PORTEN_B12 ,PORTEN_B20 ,PORTEN_B13 ,PORTEN_B21 ,PORTEN_B14 ,PORTEN_B22 ,PORTEN_B15
 ,PORTEN_B23 ,PORTEN_B16 ,PORTEN_B24 ,PORTEN_B17 ,PORTEN_B25 ,PORTEN_B18 ,PORTEN_B26 ,PORTEN_B19
);

  input CLK30MHZ ;
  input EVAOSCMCLK ;
  input RESET_B ;
  input ICESYSRES_B ;
  input ICECPURES_B ;
  input EACONNECT_B ;
  input TCCONNECT_B ;
  input TVDDON ;
  input USBCLK ;
  input USBRD_B ;
  input USBWR0_B ;
  input USBA1 ;
  input USBA2 ;
  input USBA3 ;
  input USBA4 ;
  input USBA19 ;
  input USBA20 ;
  input USBA21 ;
  input EROMPD32 ;
  input EROMPD33 ;
  input EROMPD34 ;
  input EROMPD35 ;
  input P121 ;
  input P122 ;
  input P123 ;
  input P124 ;
  input PTTL03 ;
  input PTTL11 ;
  input PTTL04 ;
  input PTTL10 ;
  input PTTL13 ;
  input PTTL14 ;
  input PTTL15 ;
  input PTTL16 ;
  input PTTL17 ;
  input P137 ;
  input ADINT_B ;
  input AD_DB9 ;
  input AD_DB8 ;
  input AD_DB7 ;
  input AD_DB6 ;
  input AD_DB5 ;
  input AD_DB4 ;
  input AD_DB3 ;
  input AD_DB2 ;
  input AD_DB1 ;
  input AD_DB0 ;

  output TVDDSEL ;
  output LEDCLOCK_B ;
  output LEDRESET_B ;
  output LEDRUN_B ;
  output LEDSTANDBY_B ;
  output LEDTVDD_B ;
  output LEDWAIT_B ;
  output USBWAIT_B ;
  output PPUP0 ;
  output PPUP1 ;
  output PPUP2 ;
  output PPUP15 ;
  output PPUP31 ;
  output PPUP4 ;
  output PPUP5 ;
  output PPUP6 ;
  output PPUP7 ;
  output PPUP8 ;
  output PPUP9 ;
  output PPUP18 ;
  output PPUP26 ;
  output PPUP19 ;
  output PPUP27 ;
  output PPUP28 ;
  output PPUP29 ;
  output EROMCLK ;
  output EROMCSB ;
  output EROMPA2 ;
  output EROMWRB ;
  output EROMRDB ;
  output EROMPA0 ;
  output EROMPA1 ;
  output EROMPA3 ;
  output EROMPA4 ;
  output EROMPA5 ;
  output EROMPA6 ;
  output EROMPA7 ;
  output EROMPA8 ;
  output EROMPA9 ;
  output EROMPA10 ;
  output EROMPA11 ;
  output EROMPA12 ;
  output EROMPA13 ;
  output EROMPA14 ;
  output EROMPA15 ;
  output EROMPA16 ;
  output EROMPA17 ;
  output DIS_OUT ;
  output WWR_OUT ;
  output MRG00_OUT ;
  output MRG01_OUT ;
  output MRG10_OUT ;
  output MRG11_OUT ;
  output MRG12_OUT ;
  output READ_OUT ;
  output FCLK_OUT ;
  output RDCLKP1_OUT ;
  output PROGI_OUT ;
  output CER_OUT ;
  output SER_OUT ;
  output EXA_OUT ;
  output EXER_OUT ;
  output BFA_OUT ;
  output TMEMCLK0 ;
  output TMEMCLK1 ;
  output TMEMCLK2 ;
  output TMEMCS_B ;
  output TMEMRD_B ;
  output TMEMWR_B ;
  output TMEMA0 ;
  output TMEMA1 ;
  output TMEMA2 ;
  output TMEMA3 ;
  output TMEMA4 ;
  output TMEMA5 ;
  output TMEMA6 ;
  output TMEMA7 ;
  output TMEMA8 ;
  output TMEMA9 ;
  output TMEMA10 ;
  output TMEMA11 ;
  output TMEMA12 ;
  output TMEMA13 ;
  output TMEMA14 ;
  output TMEMA15 ;
  output TMEMA16 ;
  output LVISEL ;
  output P130 ;
  output AP10 ;
  output AP11 ;
  output AP12 ;
  output AP20 ;
  output AP1 ;
  output AP2 ;
  output AP3 ;
  output AP4 ;
  output AP5 ;
  output AP6 ;
  output AP7 ;
  output AP8 ;
  output AP9 ;
  output AP17 ;
  output AP25 ;
  output AP33 ;
  output AP41 ;
  output AP13 ;
  output AP21 ;
  output AP18 ;
  output AP26 ;
  output AP34 ;
  output AP42 ;
  output AP50 ;
  output AP19 ;
  output AP27 ;
  output AP35 ;
  output AP43 ;
  output AP51 ;
  output PPUP3 ;
  output PPUP10 ;
  output PPUP11 ;
  output PPUP12 ;
  output PPUP20 ;
  output PPUP13 ;
  output PPUP21 ;
  output PPUP14 ;
  output PPUP30 ;
  output PPUP16 ;
  output PPUP24 ;
  output PPUP17 ;
  output PPUP25 ;
  output PUPLE0 ;
  output PUPLE1 ;
  output PUPLE2 ;
  output PUPLE3 ;
  output PUPLE4 ;
  output PUPLE5 ;
  output PSSC0 ;
  output PSSC1 ;
  output PSSC2 ;
  output PSSC3 ;
  output PSSC4 ;
  output PSSC5 ;
  output PIO00 ;
  output PIO01 ;
  output PIO02 ;
  output PIO10 ;
  output PIO03 ;
  output PIO11 ;
  output PIO04 ;
  output PIO12 ;
  output PIO20 ;
  output PIO05 ;
  output PIO13 ;
  output PIO21 ;
  output PIO06 ;
  output PIO14 ;
  output PIO22 ;
  output PIO30 ;
  output PIO15 ;
  output PIO23 ;
  output PIO31 ;
  output PIO16 ;
  output PIO24 ;
  output PIO40 ;
  output PIO17 ;
  output PIO25 ;
  output PIO41 ;
  output PIO26 ;
  output PIO42 ;
  output PIO50 ;
  output PIO27 ;
  output PIO43 ;
  output PIO51 ;
  output PIO52 ;
  output PIO60 ;
  output PIO53 ;
  output PIO61 ;
  output PIO54 ;
  output PIO62 ;
  output PIO70 ;
  output PIO55 ;
  output PIO63 ;
  output PIO71 ;
  output PIO72 ;
  output PIO73 ;
  output PIO74 ;
  output PIO75 ;
  output PIO76 ;
  output PIO77 ;
  output PIO120 ;
  output PIO121 ;
  output PIO122 ;
  output PIO130 ;
  output PIO123 ;
  output PIO124 ;
  output PIO140 ;
  output PIO141 ;
  output PIO146 ;
  output PIO147 ;
  output ADCS_B ;
  output ADRD_B ;
  output ADSH_B ;
  output AD_A4 ;
  output AD_A3 ;
  output AD_A2 ;
  output AD_A1 ;
  output AD_A0 ;
  output ADGSELMOD ;
  output PORTEN_B0 ;
  output PORTEN_B1 ;
  output PORTEN_B2 ;
  output PORTEN_B3 ;
  output PORTEN_B4 ;
  output PORTEN_B5 ;
  output PORTEN_B6 ;
  output PORTEN_B7 ;
  output PORTEN_B8 ;
  output PORTEN_B9 ;
  output PORTEN_B10 ;
  output PORTEN_B11 ;
  output EMVDDSEL_B ;
  output ADVSELMOD ;
  output AP14 ;
  output AP22 ;
  output AP30 ;
  output AP15 ;
  output AP23 ;
  output AP31 ;
  output AP16 ;
  output AP24 ;
  output AP32 ;
  output AP40 ;
  output AP28 ;
  output AP36 ;
  output AP44 ;
  output AP52 ;
  output AP60 ;
  output AP29 ;
  output AP37 ;
  output AP45 ;
  output AP53 ;
  output AP61 ;
  output AP38 ;
  output AP46 ;
  output AP54 ;
  output AP62 ;
  output AP39 ;
  output AP47 ;
  output AP55 ;
  output AP63 ;
  output AP48 ;
  output AP56 ;
  output AP64 ;
  output AP49 ;
  output AP57 ;
  output AP65 ;
  output AP58 ;
  output AP59 ;
  output APIO1 ;
  output APIO2 ;
  output APIO3 ;
  output APIO4 ;
  output APIO5 ;
  output APIO6 ;
  output APIO7 ;
  output APIO8 ;
  output APIO9 ;
  output APIO10 ;
  output APIO11 ;
  output APIO12 ;
  output APIO20 ;
  output APIO13 ;
  output APIO21 ;
  output APIO14 ;
  output APIO22 ;
  output APIO30 ;
  output APIO15 ;
  output APIO23 ;
  output APIO31 ;
  output APIO16 ;
  output APIO24 ;
  output APIO32 ;
  output APIO40 ;
  output APIO17 ;
  output APIO25 ;
  output APIO33 ;
  output APIO41 ;
  output APIO18 ;
  output APIO26 ;
  output APIO34 ;
  output APIO42 ;
  output APIO50 ;
  output APIO19 ;
  output APIO27 ;
  output APIO35 ;
  output APIO43 ;
  output APIO51 ;
  output APIO28 ;
  output APIO36 ;
  output APIO44 ;
  output APIO52 ;
  output APIO60 ;
  output APIO29 ;
  output APIO37 ;
  output APIO45 ;
  output APIO53 ;
  output APIO61 ;
  output APIO38 ;
  output APIO46 ;
  output APIO54 ;
  output APIO62 ;
  output APIO39 ;
  output APIO47 ;
  output APIO55 ;
  output APIO63 ;
  output APIO48 ;
  output APIO56 ;
  output APIO64 ;
  output APIO49 ;
  output APIO57 ;
  output APIO65 ;
  output APIO58 ;
  output APIO59 ;
  output PIO_ANALOG0 ;
  output PIO_ANALOG1 ;
  output PIO_ANALOG2 ;
  output PIO_ANALOG3 ;
  output PIO_ANALOG4 ;
  output PIO_ANALOG5 ;
  output PORTEN_B12 ;
  output PORTEN_B20 ;
  output PORTEN_B13 ;
  output PORTEN_B21 ;
  output PORTEN_B14 ;
  output PORTEN_B22 ;
  output PORTEN_B15 ;
  output PORTEN_B23 ;
  output PORTEN_B16 ;
  output PORTEN_B24 ;
  output PORTEN_B17 ;
  output PORTEN_B25 ;
  output PORTEN_B18 ;
  output PORTEN_B26 ;
  output PORTEN_B19 ;

  inout USBD0 ;
  inout USBD1 ;
  inout USBD2 ;
  inout USBD3 ;
  inout USBD4 ;
  inout USBD5 ;
  inout USBD6 ;
  inout USBD7 ;
  inout USBD8 ;
  inout USBD9 ;
  inout USBD10 ;
  inout USBD11 ;
  inout USBD12 ;
  inout USBD13 ;
  inout USBD14 ;
  inout USBD15 ;
  inout EROMPD0 ;
  inout EROMPD1 ;
  inout EROMPD2 ;
  inout EROMPD3 ;
  inout EROMPD4 ;
  inout EROMPD5 ;
  inout EROMPD6 ;
  inout EROMPD7 ;
  inout EROMPD8 ;
  inout EROMPD9 ;
  inout EROMPD10 ;
  inout EROMPD11 ;
  inout EROMPD12 ;
  inout EROMPD20 ;
  inout EROMPD13 ;
  inout EROMPD21 ;
  inout EROMPD14 ;
  inout EROMPD22 ;
  inout EROMPD30 ;
  inout EROMPD15 ;
  inout EROMPD23 ;
  inout EROMPD31 ;
  inout EROMPD16 ;
  inout EROMPD24 ;
  inout EROMPD17 ;
  inout EROMPD25 ;
  inout EROMPD18 ;
  inout EROMPD26 ;
  inout EROMPD19 ;
  inout EROMPD27 ;
  inout EROMPD28 ;
  inout EROMPD29 ;
  inout TMEMD0 ;
  inout TMEMD1 ;
  inout TMEMD2 ;
  inout TMEMD3 ;
  inout TMEMD4 ;
  inout TMEMD5 ;
  inout TMEMD6 ;
  inout TMEMD7 ;
  inout TMEMD8 ;
  inout TMEMD9 ;
  inout TMEMD10 ;
  inout TMEMD11 ;
  inout TMEMD12 ;
  inout TMEMD20 ;
  inout TMEMD13 ;
  inout TMEMD21 ;
  inout TMEMD14 ;
  inout TMEMD22 ;
  inout TMEMD30 ;
  inout TMEMD15 ;
  inout TMEMD23 ;
  inout TMEMD31 ;
  inout TMEMD16 ;
  inout TMEMD24 ;
  inout TMEMD32 ;
  inout TMEMD40 ;
  inout TMEMD17 ;
  inout TMEMD25 ;
  inout TMEMD33 ;
  inout TMEMD41 ;
  inout TMEMD18 ;
  inout TMEMD26 ;
  inout TMEMD34 ;
  inout TMEMD42 ;
  inout TMEMD50 ;
  inout TMEMD19 ;
  inout TMEMD27 ;
  inout TMEMD35 ;
  inout TMEMD43 ;
  inout TMEMD51 ;
  inout TMEMD28 ;
  inout TMEMD36 ;
  inout TMEMD44 ;
  inout TMEMD52 ;
  inout TMEMD60 ;
  inout TMEMD29 ;
  inout TMEMD37 ;
  inout TMEMD45 ;
  inout TMEMD53 ;
  inout TMEMD61 ;
  inout TMEMD38 ;
  inout TMEMD46 ;
  inout TMEMD54 ;
  inout TMEMD62 ;
  inout TMEMD70 ;
  inout TMEMD39 ;
  inout TMEMD47 ;
  inout TMEMD55 ;
  inout TMEMD63 ;
  inout TMEMD71 ;
  inout TMEMD48 ;
  inout TMEMD56 ;
  inout TMEMD64 ;
  inout TMEMD72 ;
  inout TMEMD80 ;
  inout TMEMD49 ;
  inout TMEMD57 ;
  inout TMEMD65 ;
  inout TMEMD73 ;
  inout TMEMD81 ;
  inout TMEMD58 ;
  inout TMEMD66 ;
  inout TMEMD74 ;
  inout TMEMD82 ;
  inout TMEMD90 ;
  inout TMEMD59 ;
  inout TMEMD67 ;
  inout TMEMD75 ;
  inout TMEMD83 ;
  inout TMEMD91 ;
  inout TMEMD68 ;
  inout TMEMD76 ;
  inout TMEMD84 ;
  inout TMEMD92 ;
  inout TMEMD69 ;
  inout TMEMD77 ;
  inout TMEMD85 ;
  inout TMEMD93 ;
  inout TMEMD78 ;
  inout TMEMD86 ;
  inout TMEMD94 ;
  inout TMEMD79 ;
  inout TMEMD87 ;
  inout TMEMD95 ;
  inout TMEMD88 ;
  inout TMEMD96 ;
  inout TMEMD89 ;
  inout TMEMD97 ;
  inout TMEMD98 ;
  inout TMEMD99 ;
  inout TMEMD100 ;
  inout TMEMD101 ;
  inout TMEMD102 ;
  inout TMEMD103 ;
  inout TMEMD104 ;
  inout TMEMD105 ;
  inout TMEMD106 ;
  inout TMEMD107 ;
  inout P140 ;
  inout P00 ;
  inout P01 ;
  inout P02 ;
  inout P10 ;
  inout P03 ;
  inout P11 ;
  inout P04 ;
  inout P12 ;
  inout P20 ;
  inout P05 ;
  inout P13 ;
  inout P21 ;
  inout P06 ;
  inout P14 ;
  inout P22 ;
  inout P30 ;
  inout P15 ;
  inout P23 ;
  inout P31 ;
  inout P16 ;
  inout P24 ;
  inout P40 ;
  inout P17 ;
  inout P25 ;
  inout P41 ;
  inout P26 ;
  inout P42 ;
  inout P50 ;
  inout P27 ;
  inout P43 ;
  inout P51 ;
  inout P52 ;
  inout P60 ;
  inout P53 ;
  inout P61 ;
  inout P54 ;
  inout P62 ;
  inout P70 ;
  inout P55 ;
  inout P63 ;
  inout P71 ;
  inout P72 ;
  inout P73 ;
  inout P74 ;
  inout P75 ;
  inout P76 ;
  inout P77 ;
  inout P120 ;
  inout P141 ;
  inout P146 ;
  inout P147 ;
 
  wire  CLK30MHZ ,EVAOSCMCLK ,RESET_B ,ICESYSRES_B ,ICECPURES_B ,EACONNECT_B ,TCCONNECT_B ,TVDDSEL ;
  wire  TVDDON ,LEDCLOCK_B ,LEDRESET_B ,LEDRUN_B ,LEDSTANDBY_B ,LEDTVDD_B ,LEDWAIT_B ,USBCLK ;
  wire  USBRD_B ,USBWR0_B ,USBWAIT_B ,USBA1 ,PROGI ,USBA2 ,PPUP0 ,USBA3 ;
  wire  PPUP1 ,USBA4 ,PPUP2 ,USBA19 ,PPUP15 ,PPUP31 ,USBA20 ,USBA21 ;
  wire  USBD0 ,PPUP4 ,USBD1 ,PPUP5 ,USBD2 ,PPUP6 ,USBD3 ,PPUP7 ;
  wire  USBD4 ,PPUP8 ,USBD5 ,PPUP9 ,USBD6 ,USBD7 ,USBD8 ,USBD9 ;
  wire  USBD10 ,PPUP18 ,PPUP26 ,USBD11 ,PPUP19 ,PPUP27 ,USBD12 ,PPUP28 ;
  wire  USBD13 ,PPUP29 ,USBD14 ,USBD15 ,EROMCLK ,EROMCSB ,EROMPA2 ,EROMWRB ;
  wire  EROMRDB ,EROMPA0 ,EROMPA1 ,EROMPA3 ,EROMPA4 ,EROMPA5 ,EROMPA6 ,EROMPD0 ;
  wire  EROMPA7 ,EROMPD1 ,EROMPA8 ,EROMPD2 ,EROMPA9 ,EROMPD3 ,EROMPA10 ,EROMPA11 ;
  wire  EROMPA12 ,EROMPA13 ,EROMPA14 ,EROMPA15 ,EROMPA16 ,EROMPA17 ,EROMPD4 ,EROMPD5 ;
  wire  EROMPD6 ,EROMPD7 ,EROMPD8 ,EROMPD9 ,EROMPD10 ,EROMPD11 ,EROMPD12 ,EROMPD20 ;
  wire  EROMPD13 ,EROMPD21 ,EROMPD14 ,EROMPD22 ,EROMPD30 ,EROMPD15 ,EROMPD23 ,EROMPD31 ;
  wire  EROMPD16 ,EROMPD24 ,EROMPD32 ,EROMPD17 ,EROMPD25 ,EROMPD33 ,EROMPD18 ,EROMPD26 ;
  wire  EROMPD34 ,EROMPD19 ,EROMPD27 ,EROMPD35 ,EROMPD28 ,EROMPD29 ,DIS_OUT ,WWR_OUT ;
  wire  MRG00_OUT ,MRG01_OUT ,MRG10_OUT ,MRG11_OUT ,MRG12_OUT ,READ_OUT ,FCLK_OUT ,RDCLKP1_OUT ;
  wire  PROGI_OUT ,CER_OUT ,SER_OUT ,EXA_OUT ,EXER_OUT ,BFA_OUT ,TMEMCLK0 ,TMEMCLK1 ;
  wire  TMEMCLK2 ,TMEMCS_B ,TMEMRD_B ,TMEMWR_B ,TMEMA0 ,TMEMA1 ,TMEMA2 ,TMEMA3 ;
  wire  TMEMA4 ,TMEMA5 ,TMEMA6 ,TMEMD0 ,TMEMA7 ,TMEMD1 ,TMEMA8 ,TMEMD2 ;
  wire  TMEMA9 ,TMEMD3 ,TMEMA10 ,TMEMA11 ,TMEMA12 ,TMEMA13 ,TMEMA14 ,SLFLASH ;
  wire  WAITFL2 ,TMEMA15 ,TMEMA16 ,TMEMD4 ,TMEMD5 ,TMEMD6 ,TMEMD7 ,TMEMD8 ;
  wire  TMEMD9 ,TMEMD10 ,TMEMD11 ,TMEMD12 ,TMEMD20 ,TMEMD13 ,TMEMD21 ,TMEMD14 ;
  wire  TMEMD22 ,TMEMD30 ,TMEMD15 ,TMEMD23 ,TMEMD31 ,TMEMD16 ,TMEMD24 ,TMEMD32 ;
  wire  TMEMD40 ,TMEMD17 ,TMEMD25 ,TMEMD33 ,TMEMD41 ,TMEMD18 ,TMEMD26 ,TMEMD34 ;
  wire  TMEMD42 ,TMEMD50 ,TMEMD19 ,TMEMD27 ,TMEMD35 ,TMEMD43 ,TMEMD51 ,TMEMD28 ;
  wire  TMEMD36 ,TMEMD44 ,TMEMD52 ,TMEMD60 ,TMEMD29 ,TMEMD37 ,TMEMD45 ,TMEMD53 ;
  wire  TMEMD61 ,TMEMD38 ,TMEMD46 ,TMEMD54 ,TMEMD62 ,TMEMD70 ,TMEMD39 ,TMEMD47 ;
  wire  TMEMD55 ,TMEMD63 ,TMEMD71 ,TMEMD48 ,TMEMD56 ,TMEMD64 ,TMEMD72 ,TMEMD80 ;
  wire  TMEMD49 ,TMEMD57 ,TMEMD65 ,TMEMD73 ,TMEMD81 ,TMEMD58 ,TMEMD66 ,TMEMD74 ;
  wire  TMEMD82 ,TMEMD90 ,TMEMD59 ,TMEMD67 ,TMEMD75 ,TMEMD83 ,TMEMD91 ,TMEMD68 ;
  wire  TMEMD76 ,TMEMD84 ,TMEMD92 ,TMEMD69 ,TMEMD77 ,TMEMD85 ,TMEMD93 ,TMEMD78 ;
  wire  TMEMD86 ,TMEMD94 ,TMEMD79 ,TMEMD87 ,TMEMD95 ,TMEMD88 ,TMEMD96 ,TMEMD89 ;
  wire  TMEMD97 ,TMEMD98 ,TMEMD99 ,TMEMD100 ,TMEMD101 ,TMEMD102 ,TMEMD103 ,TMEMD104 ;
  wire  TMEMD105 ,TMEMD106 ,TMEMD107 ,LVISEL ,PREFIX ,P121 ,P122 ,P130 ;
  wire  AP10 ,P123 ,AP11 ,P124 ,P140 ,AP12 ,AP20 ,P00 ;
  wire  P01 ,P02 ,P10 ,P03 ,P11 ,PTTL03 ,PTTL11 ,P04 ;
  wire  P12 ,P20 ,PTTL04 ,P05 ,P13 ,P21 ,AP1 ,BFA ;
  wire  P06 ,P14 ,P22 ,P30 ,AP2 ,PTTL10 ,PTTL13 ,PTTL14 ;
  wire  P15 ,P23 ,P31 ,AP3 ,PTTL15 ,P16 ,P24 ,P40 ;
  wire  AP4 ,PTTL16 ,P17 ,P25 ,P41 ,AP5 ,PTTL17 ,P26 ;
  wire  P42 ,P50 ,AP6 ,P27 ,P43 ,P51 ,AP7 ,P52 ;
  wire  P60 ,AP8 ,P53 ,P61 ,AP9 ,P54 ,P62 ,P70 ;
  wire  P55 ,P63 ,P71 ,P72 ,P73 ,P74 ,P75 ,P76 ;
  wire  P77 ,P120 ,P137 ,AP17 ,AP25 ,AP33 ,AP41 ,P141 ;
  wire  AP13 ,AP21 ,P146 ,AP18 ,AP26 ,AP34 ,AP42 ,AP50 ;
  wire  P147 ,AP19 ,AP27 ,AP35 ,AP43 ,AP51 ,PPUP3 ,PPUP10 ;
  wire  PPUP11 ,PPUP12 ,PPUP20 ,PPUP13 ,PPUP21 ,PPUP14 ,PPUP30 ,PPUP16 ;
  wire  PPUP24 ,PPUP17 ,PPUP25 ,PUPLE0 ,PUPLE1 ,PUPLE2 ,PUPLE3 ,PUPLE4 ;
  wire  PUPLE5 ,PSSC0 ,PSSC1 ,SLMEM ,PSSC2 ,PSSC3 ,PSSC4 ,PSSC5 ;
  wire  PIO00 ,PIO01 ,PIO02 ,PIO10 ,PIO03 ,PIO11 ,PIO04 ,PIO12 ;
  wire  PIO20 ,PIO05 ,PIO13 ,PIO21 ,PIO06 ,PIO14 ,PIO22 ,PIO30 ;
  wire  PIO15 ,PIO23 ,PIO31 ,PIO16 ,PIO24 ,PIO40 ,PIO17 ,PIO25 ;
  wire  PIO41 ,PIO26 ,PIO42 ,PIO50 ,PIO27 ,PIO43 ,PIO51 ,PIO52 ;
  wire  PIO60 ,PIO53 ,PIO61 ,PIO54 ,PIO62 ,PIO70 ,PIO55 ,PIO63 ;
  wire  PIO71 ,PIO72 ,PIO73 ,PIO74 ,PIO75 ,PIO76 ,PIO77 ,PIO120 ;
  wire  PIO121 ,PIO122 ,PIO130 ,PIO123 ,PIO124 ,PIO140 ,PIO141 ,PIO146 ;
  wire  PIO147 ,ADINT_B ,P05PUON ,P13PUON ,AD_DB9 ,AD_DB8 ,AD_DB7 ,AD_DB6 ;
  wire  AD_DB5 ,P77ENI ,AD_DB4 ,AD_DB3 ,P76ENO ,AD_DB2 ,AD_DB1 ,AD_DB0 ;
  wire  ADCS_B ,ADRD_B ,P74DIN ,ADSH_B ,P77DIN ,AD_A4 ,AD_A3 ,AD_A2 ;
  wire  AD_A1 ,AD_A0 ,ADGSELMOD ,PORTEN_B0 ,PORTEN_B1 ,PORTEN_B2 ,PORTEN_B3 ,PORTEN_B4 ;
  wire  PORTEN_B5 ,PORTEN_B6 ,PORTEN_B7 ,PORTEN_B8 ,PORTEN_B9 ,PORTEN_B10 ,PORTEN_B11 ,EMVDDSEL_B ;
  wire  ADVSELMOD ,AP14 ,AP22 ,AP30 ,AP15 ,AP23 ,AP31 ,AP16 ;
  wire  AP24 ,AP32 ,AP40 ,AP28 ,AP36 ,AP44 ,AP52 ,AP60 ;
  wire  AP29 ,AP37 ,AP45 ,AP53 ,AP61 ,AP38 ,AP46 ,AP54 ;
  wire  AP62 ,DCE0 ,AP39 ,AP47 ,AP55 ,AP63 ,AP48 ,AP56 ;
  wire  AP64 ,AP49 ,AP57 ,AP65 ,AP58 ,AP59 ,APIO1 ,APIO2 ;
  wire  APIO3 ,APIO4 ,APIO5 ,APIO6 ,APIO7 ,APIO8 ,APIO9 ,APIO10 ;
  wire  APIO11 ,APIO12 ,APIO20 ,APIO13 ,APIO21 ,APIO14 ,APIO22 ,APIO30 ;
  wire  APIO15 ,APIO23 ,APIO31 ,APIO16 ,APIO24 ,APIO32 ,APIO40 ,APIO17 ;
  wire  APIO25 ,APIO33 ,APIO41 ,APIO18 ,APIO26 ,APIO34 ,APIO42 ,APIO50 ;
  wire  APIO19 ,APIO27 ,APIO35 ,APIO43 ,APIO51 ,APIO28 ,APIO36 ,APIO44 ;
  wire  APIO52 ,APIO60 ,APIO29 ,APIO37 ,APIO45 ,APIO53 ,APIO61 ,APIO38 ;
  wire  APIO46 ,APIO54 ,APIO62 ,APIO39 ,APIO47 ,APIO55 ,APIO63 ,APIO48 ;
  wire  APIO56 ,APIO64 ,APIO49 ,APIO57 ,APIO65 ,APIO58 ,APIO59 ,FCHRAM ;
  wire  PIO_ANALOG0 ,PIO_ANALOG1 ,PIO_ANALOG2 ,PIO_ANALOG3 ,PIO_ANALOG4 ,PIO_ANALOG5 ,PORTEN_B12 ,PORTEN_B20 ;
  wire  PORTEN_B13 ,PORTEN_B21 ,PORTEN_B14 ,PORTEN_B22 ,PORTEN_B15 ,PORTEN_B23 ,PORTEN_B16 ,PORTEN_B24 ;
  wire  PORTEN_B17 ,PORTEN_B25 ,PORTEN_B18 ,PORTEN_B26 ,PORTEN_B19 ,FCLK_ICE ,PSEUDOON2 ,PSEUDOON3 ;
  wire  PSEUDOON4 ,PSEUDOON5 ,PSEUDOON6 ,PSEUDOON7 ,FCLK1 ,FLSPM ,RO137 ,RO129 ;
  wire  EXMA3 ,DRO00 ,DRO01 ,DRO02 ,DRO03 ,DRO04 ,DRO05 ,DRO06 ;
  wire  DRO07 ,DRO08 ,DRO09 ,DRO010 ,DRO011 ,ICEMKLVI ,ICEMKWDT ,RESINB ;
  wire  RESETB ,SBANDOCD ,LOCK64FAIL ,LOCK48FAIL ,LOCKHROSCFAIL ,SYSRSOUTB ,P30PUONOUT ,P14PUONOUT ;
  wire  P06PUONOUT ,P31PUONOUT ,P15PUONOUT ,P70PUONOUT ,P54PUONOUT ,P71PUONOUT ,P55PUONOUT ,P72PUONOUT ;
  wire  P73PUONOUT ,P74PUONOUT ,P75PUONOUT ,P76PUONOUT ,P77PUONOUT ,P10PUONOUT ,P02PUONOUT ,P11PUONOUT ;
  wire  P03PUONOUT ,P12PUONOUT ,P04PUONOUT ,P13PUONOUT ,P05PUONOUT ,P16PUONOUT ,P40PUONOUT ,P17PUONOUT ;
  wire  P41PUONOUT ,P42PUONOUT ,P50PUONOUT ,P43PUONOUT ,P51PUONOUT ,P52PUONOUT ,P53PUONOUT ,P00PUONOUT ;
  wire  P01PUONOUT ,P140PUONOUT ,P141PUONOUT ,P146PUONOUT ,P120PUONOUT ,P147PUONOUT ,pull_down0 ,pull_down1 ;
  wire  pull_down2 ,pull_down3 ,pull_down4 ,pull_down5 ,pull_down6 ,pull_down7 ,pull_down8 ,pull_down9 ;
  wire  pull_down10 ,pull_down11 ,pull_down12 ,pull_down20 ,pull_down13 ,pull_down21 ,pull_down14 ,pull_down22 ;
  wire  pull_down30 ,pull_down15 ,pull_down23 ,pull_down31 ,pull_down16 ,pull_down24 ,pull_down32 ,pull_down40 ;
  wire  pull_down17 ,pull_down25 ,pull_down33 ,pull_down41 ,pull_down18 ,pull_down26 ,pull_down34 ,pull_down42 ;
  wire  pull_down50 ,pull_down19 ,pull_down27 ,pull_down35 ,pull_down43 ,pull_down51 ,pull_down28 ,pull_down36 ;
  wire  pull_down44 ,pull_down52 ,pull_down60 ,pull_down29 ,pull_down37 ,pull_down45 ,pull_down53 ,pull_down61 ;
  wire  pull_down38 ,pull_down46 ,pull_down54 ,pull_down62 ,pull_down70 ,pull_down39 ,pull_down47 ,pull_down55 ;
  wire  pull_down63 ,pull_down71 ,pull_down48 ,pull_down56 ,pull_down64 ,pull_down72 ,pull_down80 ,pull_down49 ;
  wire  pull_down57 ,pull_down65 ,pull_down73 ,pull_down81 ,pull_down58 ,pull_down66 ,pull_down74 ,pull_down82 ;
  wire  pull_down90 ,pull_down59 ,pull_down67 ,pull_down75 ,pull_down83 ,pull_down91 ,pull_down68 ,pull_down76 ;
  wire  pull_down84 ,pull_down92 ,pull_down69 ,pull_down77 ,pull_down85 ,pull_down93 ,pull_down78 ,pull_down86 ;
  wire  pull_down94 ,pull_down79 ,pull_down87 ,pull_down95 ,pull_down88 ,pull_down96 ,pull_down89 ,pull_down97 ;
  wire  pull_down98 ,pull_down99 ,pull_down100 ,pull_down101 ,pull_down102 ,pull_down110 ,pull_down103 ,pull_down111 ;
  wire  pull_down104 ,pull_down112 ,pull_down120 ,pull_down200 ,pull_down105 ,pull_down113 ,pull_down121 ,pull_down201 ;
  wire  pull_down106 ,pull_down114 ,pull_down122 ,pull_down130 ,pull_down202 ,pull_down210 ,pull_down107 ,pull_down115 ;
  wire  pull_down123 ,pull_down131 ,pull_down203 ,pull_down211 ,pull_down108 ,pull_down116 ,pull_down124 ,pull_down132 ;
  wire  pull_down140 ,pull_down204 ,pull_down212 ,pull_down220 ,pull_down300 ,pull_down109 ,pull_down117 ,pull_down125 ;
  wire  pull_down133 ,pull_down141 ,pull_down205 ,pull_down213 ,pull_down221 ,pull_down301 ,pull_down118 ,pull_down126 ;
  wire  pull_down134 ,pull_down142 ,pull_down150 ,pull_down206 ,pull_down214 ,pull_down222 ,pull_down230 ,pull_down302 ;
  wire  pull_down310 ,pull_down119 ,pull_down127 ,pull_down135 ,pull_down143 ,pull_down151 ,pull_down207 ,pull_down215 ;
  wire  pull_down223 ,pull_down231 ,pull_down303 ,pull_down311 ,pull_down128 ,pull_down136 ,pull_down144 ,pull_down152 ;
  wire  pull_down160 ,pull_down208 ,pull_down216 ,pull_down224 ,pull_down232 ,pull_down240 ,pull_down304 ,pull_down312 ;
  wire  pull_down320 ,pull_down400 ,pull_down129 ,pull_down137 ,pull_down145 ,pull_down153 ,pull_down161 ,pull_down209 ;
  wire  pull_down217 ,pull_down225 ,pull_down233 ,pull_down241 ,pull_down305 ,pull_down313 ,pull_down321 ,pull_down401 ;
  wire  pull_down138 ,pull_down146 ,pull_down154 ,pull_down162 ,pull_down170 ,pull_down218 ,pull_down226 ,pull_down234 ;
  wire  pull_down242 ,pull_down250 ,pull_down306 ,pull_down314 ,pull_down322 ,pull_down330 ,pull_down402 ,pull_down410 ;
  wire  pull_down139 ,pull_down147 ,pull_down155 ,pull_down163 ,pull_down171 ,pull_down219 ,pull_down227 ,pull_down235 ;
  wire  pull_down243 ,pull_down251 ,pull_down307 ,pull_down315 ,pull_down323 ,pull_down331 ,pull_down403 ,pull_down411 ;
  wire  pull_down148 ,pull_down156 ,pull_down164 ,pull_down172 ,pull_down180 ,pull_down228 ,pull_down236 ,pull_down244 ;
  wire  pull_down252 ,pull_down260 ,pull_down308 ,pull_down316 ,pull_down324 ,pull_down332 ,pull_down340 ,pull_down404 ;
  wire  pull_down412 ,pull_down420 ,pull_down500 ,pull_down149 ,pull_down157 ,pull_down165 ,pull_down173 ,pull_down181 ;
  wire  pull_down229 ,pull_down237 ,pull_down245 ,pull_down253 ,pull_down261 ,pull_down309 ,pull_down317 ,pull_down325 ;
  wire  pull_down333 ,pull_down341 ,pull_down405 ,pull_down413 ,pull_down421 ,pull_down501 ,pull_down158 ,pull_down166 ;
  wire  pull_down174 ,pull_down182 ,pull_down190 ,pull_down238 ,pull_down246 ,pull_down254 ,pull_down262 ,pull_down270 ;
  wire  pull_down318 ,pull_down326 ,pull_down334 ,pull_down342 ,pull_down350 ,pull_down406 ,pull_down414 ,pull_down422 ;
  wire  pull_down430 ,pull_down502 ,pull_down510 ,pull_down159 ,pull_down167 ,pull_down175 ,pull_down183 ,pull_down191 ;
  wire  pull_down239 ,pull_down247 ,pull_down255 ,pull_down263 ,pull_down271 ,pull_down319 ,pull_down327 ,pull_down335 ;
  wire  pull_down343 ,pull_down351 ,pull_down407 ,pull_down415 ,pull_down423 ,pull_down431 ,pull_down503 ,pull_down511 ;
  wire  pull_down168 ,pull_down176 ,pull_down184 ,pull_down192 ,pull_down248 ,pull_down256 ,pull_down264 ,pull_down272 ;
  wire  pull_down280 ,pull_down328 ,pull_down336 ,pull_down344 ,pull_down352 ,pull_down360 ,pull_down408 ,pull_down416 ;
  wire  pull_down424 ,pull_down432 ,pull_down440 ,pull_down504 ,pull_down512 ,pull_down520 ,pull_down600 ,pull_down169 ;
  wire  pull_down177 ,pull_down185 ,pull_down193 ,pull_down249 ,pull_down257 ,pull_down265 ,pull_down273 ,pull_down281 ;
  wire  pull_down329 ,pull_down337 ,pull_down345 ,pull_down353 ,pull_down361 ,pull_down409 ,pull_down417 ,pull_down425 ;
  wire  pull_down433 ,pull_down441 ,pull_down505 ,pull_down513 ,pull_down521 ,pull_down601 ,pull_down178 ,pull_down186 ;
  wire  pull_down194 ,pull_down258 ,pull_down266 ,pull_down274 ,pull_down282 ,pull_down290 ,pull_down338 ,pull_down346 ;
  wire  pull_down354 ,pull_down362 ,pull_down370 ,pull_down418 ,pull_down426 ,pull_down434 ,pull_down442 ,pull_down450 ;
  wire  pull_down506 ,pull_down514 ,pull_down522 ,pull_down530 ,pull_down602 ,pull_down610 ,pull_down179 ,pull_down187 ;
  wire  pull_down195 ,pull_down259 ,pull_down267 ,pull_down275 ,pull_down283 ,pull_down291 ,pull_down339 ,pull_down347 ;
  wire  pull_down355 ,pull_down363 ,pull_down371 ,pull_down419 ,pull_down427 ,pull_down435 ,pull_down443 ,pull_down451 ;
  wire  pull_down507 ,pull_down515 ,pull_down523 ,pull_down531 ,pull_down603 ,pull_down611 ,pull_down188 ,pull_down196 ;
  wire  pull_down268 ,pull_down276 ,pull_down284 ,pull_down292 ,pull_down348 ,pull_down356 ,pull_down364 ,pull_down372 ;
  wire  pull_down380 ,pull_down428 ,pull_down436 ,pull_down444 ,pull_down452 ,pull_down460 ,pull_down508 ,pull_down516 ;
  wire  pull_down524 ,pull_down532 ,pull_down540 ,pull_down604 ,pull_down612 ,pull_down620 ,pull_down700 ,pull_down189 ;
  wire  pull_down197 ,pull_down269 ,pull_down277 ,pull_down285 ,pull_down293 ,pull_down349 ,pull_down357 ,pull_down365 ;
  wire  pull_down373 ,pull_down381 ,pull_down429 ,pull_down437 ,pull_down445 ,pull_down453 ,pull_down461 ,pull_down509 ;
  wire  pull_down517 ,pull_down525 ,pull_down533 ,pull_down541 ,pull_down605 ,pull_down613 ,pull_down621 ,pull_down701 ;
  wire  pull_down198 ,pull_down278 ,pull_down286 ,pull_down294 ,pull_down358 ,pull_down366 ,pull_down374 ,pull_down382 ;
  wire  pull_down390 ,pull_down438 ,pull_down446 ,pull_down454 ,pull_down462 ,pull_down470 ,pull_down518 ,pull_down526 ;
  wire  pull_down534 ,pull_down542 ,pull_down550 ,pull_down606 ,pull_down614 ,pull_down622 ,pull_down630 ,pull_down702 ;
  wire  pull_down710 ,pull_down199 ,pull_down279 ,pull_down287 ,pull_down295 ,pull_down359 ,pull_down367 ,pull_down375 ;
  wire  pull_down383 ,pull_down391 ,pull_down439 ,pull_down447 ,pull_down455 ,pull_down463 ,pull_down471 ,pull_down519 ;
  wire  pull_down527 ,pull_down535 ,pull_down543 ,pull_down551 ,pull_down607 ,pull_down615 ,pull_down623 ,pull_down631 ;
  wire  pull_down703 ,pull_down711 ,pull_down288 ,pull_down296 ,pull_down368 ,pull_down376 ,pull_down384 ,pull_down392 ;
  wire  pull_down448 ,pull_down456 ,pull_down464 ,pull_down472 ,pull_down480 ,pull_down528 ,pull_down536 ,pull_down544 ;
  wire  pull_down552 ,pull_down560 ,pull_down608 ,pull_down616 ,pull_down624 ,pull_down632 ,pull_down640 ,pull_down704 ;
  wire  pull_down712 ,pull_down720 ,pull_down289 ,pull_down297 ,pull_down369 ,pull_down377 ,pull_down385 ,pull_down393 ;
  wire  pull_down449 ,pull_down457 ,pull_down465 ,pull_down473 ,pull_down481 ,pull_down529 ,pull_down537 ,pull_down545 ;
  wire  pull_down553 ,pull_down561 ,pull_down609 ,pull_down617 ,pull_down625 ,pull_down633 ,pull_down641 ,pull_down705 ;
  wire  pull_down713 ,pull_down721 ,pull_down298 ,pull_down378 ,pull_down386 ,pull_down394 ,pull_down458 ,pull_down466 ;
  wire  pull_down474 ,pull_down482 ,pull_down490 ,pull_down538 ,pull_down546 ,pull_down554 ,pull_down562 ,pull_down570 ;
  wire  pull_down618 ,pull_down626 ,pull_down634 ,pull_down642 ,pull_down650 ,pull_down706 ,pull_down714 ,pull_down722 ;
  wire  pull_down730 ,pull_down299 ,pull_down379 ,pull_down387 ,pull_down395 ,pull_down459 ,pull_down467 ,pull_down475 ;
  wire  pull_down483 ,pull_down491 ,pull_down539 ,pull_down547 ,pull_down555 ,pull_down563 ,pull_down571 ,pull_down619 ;
  wire  pull_down627 ,pull_down635 ,pull_down643 ,pull_down651 ,pull_down707 ,pull_down715 ,pull_down723 ,pull_down731 ;
  wire  pull_down388 ,pull_down396 ,pull_down468 ,pull_down476 ,pull_down484 ,pull_down492 ,pull_down548 ,pull_down556 ;
  wire  pull_down564 ,pull_down572 ,pull_down580 ,pull_down628 ,pull_down636 ,pull_down644 ,pull_down652 ,pull_down660 ;
  wire  pull_down708 ,pull_down716 ,pull_down724 ,pull_down732 ,pull_down740 ,pull_down389 ,pull_down397 ,pull_down469 ;
  wire  pull_down477 ,pull_down485 ,pull_down493 ,pull_down549 ,pull_down557 ,pull_down565 ,pull_down573 ,pull_down581 ;
  wire  pull_down629 ,pull_down637 ,pull_down645 ,pull_down653 ,pull_down661 ,pull_down709 ,pull_down717 ,pull_down725 ;
  wire  pull_down733 ,pull_down741 ,pull_down398 ,pull_down478 ,pull_down486 ,pull_down494 ,pull_down558 ,pull_down566 ;
  wire  pull_down574 ,pull_down582 ,pull_down590 ,pull_down638 ,pull_down646 ,pull_down654 ,pull_down662 ,pull_down670 ;
  wire  pull_down718 ,pull_down726 ,pull_down734 ,pull_down742 ,pull_down399 ,pull_down479 ,pull_down487 ,pull_down495 ;
  wire  pull_down559 ,pull_down567 ,pull_down575 ,pull_down583 ,pull_down591 ,pull_down639 ,pull_down647 ,pull_down655 ;
  wire  pull_down663 ,pull_down671 ,pull_down719 ,pull_down727 ,pull_down735 ,pull_down743 ,pull_down488 ,pull_down496 ;
  wire  pull_down568 ,pull_down576 ,pull_down584 ,pull_down592 ,pull_down648 ,pull_down656 ,pull_down664 ,pull_down672 ;
  wire  pull_down680 ,pull_down728 ,pull_down736 ,pull_down744 ,pull_down489 ,pull_down497 ,pull_down569 ,pull_down577 ;
  wire  pull_down585 ,pull_down593 ,pull_down649 ,pull_down657 ,pull_down665 ,pull_down673 ,pull_down681 ,pull_down729 ;
  wire  pull_down737 ,pull_down745 ,pull_down498 ,pull_down578 ,pull_down586 ,pull_down594 ,pull_down658 ,pull_down666 ;
  wire  pull_down674 ,pull_down682 ,pull_down690 ,pull_down738 ,pull_down746 ,pull_down499 ,pull_down579 ,pull_down587 ;
  wire  pull_down595 ,pull_down659 ,pull_down667 ,pull_down675 ,pull_down683 ,pull_down691 ,pull_down739 ,pull_down747 ;
  wire  pull_down588 ,pull_down596 ,pull_down668 ,pull_down676 ,pull_down684 ,pull_down692 ,pull_down589 ,pull_down597 ;
  wire  pull_down669 ,pull_down677 ,pull_down685 ,pull_down693 ,pull_down598 ,pull_down678 ,pull_down686 ,pull_down694 ;
  wire  pull_down599 ,pull_down679 ,pull_down687 ,pull_down695 ,pull_down688 ,pull_down696 ,pull_down689 ,pull_down697 ;
  wire  pull_down698 ,pull_down699 ,pull_up0 ,pull_up1 ,pull_up2 ,pull_up3 ,pull_up4 ,CIBPID31 ;
  wire  CIBPID23 ,CIBPID15 ,CIBPID30 ,CIBPID22 ,CIBPID14 ,CIBPID29 ,CIBPID28 ,CIBPID27 ;
  wire  CIBPID19 ,CIBPID26 ,CIBPID18 ,CIBPID25 ,CIBPID17 ,CIBPID24 ,CIBPID16 ,CIBPID21 ;
  wire  CIBPID13 ,CIBPID20 ,CIBPID12 ,CIBPID11 ,CIBPID10 ,CIBPID9 ,CIBPID8 ,CIBPID7 ;
  wire  CIBPID6 ,CIBPID5 ,CIBPID4 ,P42PUON ,P50PUON ,CIBPID3 ,CIBPID2 ,CIBPID1 ;
  wire  CIBPID0 ,MDRRAM15 ,MDRRAM14 ,MDRRAM13 ,MDRRAM12 ,MDRRAM11 ,MDRRAM10 ,MDRRAM9 ;
  wire  MDRRAM8 ,MDRRAM7 ,MDRRAM6 ,MDRRAM5 ,MDRRAM4 ,MDRRAM3 ,MDRRAM2 ,MDRRAM1 ;
  wire  MDRRAM0 ,ICEDO29 ,ICEDO28 ,ICEDO27 ,ICEDO19 ,ICEDO26 ,ICEDO18 ,ICEDO9 ;
  wire  ICEDO8 ,ICEDO7 ,ICEDO6 ,ICEDO5 ,ICEDO4 ,ICEDO31 ,ICEDO23 ,ICEDO15 ;
  wire  ICEDO30 ,ICEDO22 ,ICEDO14 ,ICEDO25 ,ICEDO17 ,ICEDO24 ,ICEDO16 ,ICEDO21 ;
  wire  ICEDO13 ,ICEDO20 ,ICEDO12 ,P74PUON ,ICEDO11 ,ICEDO10 ,ICEDO3 ,ICEDO2 ;
  wire  ICEDO1 ,ICEDO0 ,A19 ,A18 ,A17 ,A16 ,A15 ,A14 ;
  wire  A13 ,A12 ,A11 ,A10 ,A9 ,A8 ,A7 ,A6 ;
  wire  A5 ,A4 ,A3 ,A2 ,CE0 ,DA4 ,AF6 ,CE1 ;
  wire  DA5 ,AF7 ,SELRO1 ,CLKSEL1 ,EXA ,ICETMSPMD ,ICETMBTSEL ,BRSAM ;
  wire  RO111 ,RO031 ,RO023 ,RO015 ,RO110 ,RO030 ,RO022 ,RO014 ;
  wire  RO133 ,RO125 ,RO117 ,RO037 ,RO029 ,RO132 ,RO124 ,RO116 ;
  wire  RO036 ,RO028 ,RO131 ,RO123 ,RO115 ,RO035 ,RO027 ,RO019 ;
  wire  RO130 ,RO122 ,RO114 ,RO034 ,RO026 ,RO018 ,RO121 ,RO113 ;
  wire  RO033 ,RO025 ,RO017 ,RO120 ,RO112 ,RO032 ,RO024 ,RO016 ;
  wire  RO021 ,RO013 ,RO020 ,RO012 ,CPURD ,RO011 ,RO010 ,RO17 ;
  wire  RO09 ,RO16 ,RO08 ,RO15 ,RO07 ,RO14 ,RO06 ,RO13 ;
  wire  RO05 ,RO12 ,RO04 ,RO11 ,RO03 ,MDW9 ,RO10 ,RO02 ;
  wire  MDW8 ,RO01 ,MDW7 ,RO00 ,MDW6 ,RO136 ,RO128 ,EXMA2 ;
  wire  RO135 ,RO127 ,RO119 ,EXMA1 ,RO134 ,RO126 ,RO118 ,EXMA0 ;
  wire  RO19 ,RO18 ,DCLKSEL1 ,DRDCLKC1 ,DA13 ,AF17 ,DA12 ,AF16 ;
  wire  DA11 ,AF15 ,DA10 ,AF14 ,DA9 ,DA8 ,DA7 ,AF9 ;
  wire  DA6 ,AF8 ,DA3 ,AF5 ,DA2 ,AF4 ,DA1 ,AF3 ;
  wire  DA0 ,AF2 ,SVI ,SVVCOUT7 ,SVVCOUT6 ,SVVCOUT5 ,SVVCOUT4 ,SVVCOUT3 ;
  wire  SVVCOUT2 ,SVVCOUT1 ,SVVCOUT0 ,SVINTACK ,SOFTBRK ,ICEMSKNMI ,ICEMSKDBG ,STAGEADR1 ;
  wire  STAGEADR0 ,SKIPEXE ,PCWAITF ,CPUMASK ,CPUPID1 ,CPUMISAL ,FLREAD ,IMDR10 ;
  wire  FLREADB3 ,FLREADB2 ,FLREADB1 ,FLREADB0 ,SLEXM ,SLBMEM ,SPDEC ,SPINC ;
  wire  SPREL ,IDPOP ,MDW10 ,IMDR2 ,CPUWR ,WDOP ,ICEWAITMEM ,DMAACK ;
  wire  HLTST ,STPST ,INTACK ,OCDWAIT ,SVMOD ,SVMODF ,ALT1 ,DW21 ;
  wire  DW13 ,DRDCLK ,SLDFLASH ,ICECSGREGU ,ICEIFA4 ,ICEIFA3 ,ICEIFA2 ,PA19 ;
  wire  PC11 ,PA18 ,PC10 ,PA17 ,PA16 ,PA15 ,PA14 ,PA13 ;
  wire  DW37 ,DW29 ,PA12 ,DW36 ,DW28 ,PA11 ,DW35 ,DW27 ;
  wire  DW19 ,PA10 ,DW34 ,DW26 ,DW18 ,PA9 ,PC5 ,PA8 ;
  wire  PC4 ,PA7 ,PC3 ,PA6 ,PC2 ,PA5 ,PC1 ,DW9 ;
  wire  PA4 ,PC0 ,DW8 ,PA3 ,DW7 ,DIS ,PA2 ,DW6 ;
  wire  PC19 ,PC18 ,PC17 ,PC16 ,PC15 ,PC14 ,PC13 ,PC12 ;
  wire  PC9 ,PC8 ,PC7 ,PC6 ,IDADR31 ,IDADR23 ,IDADR15 ,ICEDI19 ;
  wire  ICEDI27 ,IDADR30 ,IDADR22 ,IDADR14 ,ICEDI18 ,ICEDI26 ,IDADR29 ,IDADR28 ;
  wire  IDADR27 ,IDADR19 ,IDADR26 ,IDADR18 ,IDADR25 ,IDADR17 ,ICEDI29 ,IDADR24 ;
  wire  IDADR16 ,ICEDI28 ,P73PUON ,IDADR21 ,IDADR13 ,ICEDI17 ,ICEDI25 ,IDADR20 ;
  wire  IDADR12 ,ICEDI16 ,ICEDI24 ,IDADR11 ,ICEDI15 ,ICEDI23 ,ICEDI31 ,IDADR10 ;
  wire  ICEDI14 ,ICEDI22 ,ICEDI30 ,IDADR9 ,IDADR8 ,IDADR7 ,ICEDI9 ,IDADR6 ;
  wire  ICEDI8 ,IDADR5 ,ICEDI7 ,IDADR4 ,ICEDI6 ,IDADR3 ,ICEDI5 ,IDADR2 ;
  wire  ICEDI4 ,IDADR1 ,ICEDI3 ,IDADR0 ,ICEDI2 ,MA15 ,MA14 ,MA13 ;
  wire  MA12 ,BEU2 ,MA11 ,BEU1 ,MA10 ,BEU0 ,MA9 ,DW1 ;
  wire  MA8 ,DW0 ,MA7 ,MA6 ,MA5 ,MA4 ,MA3 ,MA2 ;
  wire  CER ,MA1 ,MA0 ,MDW15 ,IMDR7 ,MDW14 ,IMDR6 ,MDW13 ;
  wire  IMDR5 ,MDW12 ,IMDR4 ,MDW11 ,IMDR3 ,MDW5 ,MDW4 ,MDW3 ;
  wire  MDW2 ,MDW1 ,MDW0 ,EXCH ,IMDR15 ,IMDR14 ,IMDR13 ,IMDR12 ;
  wire  IMDR11 ,IMDR9 ,IMDR8 ,IMDR1 ,IMDR0 ,CPUPID31 ,CPUPID23 ,CPUPID15 ;
  wire  CPUPID30 ,CPUPID22 ,CPUPID14 ,CPUPID29 ,CPUPID28 ,CPUPID27 ,CPUPID19 ,CPUPID26 ;
  wire  CPUPID18 ,CPUPID25 ,CPUPID17 ,CPUPID24 ,CPUPID16 ,CPUPID21 ,CPUPID13 ,CPUPID20 ;
  wire  CPUPID12 ,CPUPID11 ,CPUPID10 ,CPUPID9 ,CPUPID8 ,CPUPID7 ,CPUPID6 ,CPUPID5 ;
  wire  CPUPID4 ,CPUPID3 ,CPUPID2 ,CPUPID0 ,FLSIZE3 ,FLSIZE2 ,FLSIZE1 ,FLSIZE0 ;
  wire  RAMSIZE7 ,RAMSIZE6 ,RAMSIZE5 ,RAMSIZE4 ,RAMSIZE3 ,RAMSIZE2 ,RAMSIZE1 ,RAMSIZE0 ;
  wire  BFSIZE3 ,BFSIZE2 ,BFSIZE1 ,BFSIZE0 ,BMSIZE3 ,BMSIZE2 ,BMSIZE1 ,BMSIZE0 ;
  wire  DFSIZE1 ,DFSIZE0 ,RESB ,FCLK2 ,DW33 ,DW25 ,DW17 ,DDIS ;
  wire  DW32 ,DW24 ,DW16 ,DW31 ,DW23 ,DW15 ,DW30 ,DW22 ;
  wire  DW14 ,DW20 ,DW12 ,DW11 ,DW10 ,DW5 ,DW4 ,DW3 ;
  wire  DW2 ,TMSPMD ,TMBTSEL ,BTFLG ,READ ,RDCLKP1 ,SER ,WED ;
  wire  WWR ,MRG00 ,MRG01 ,MRG10 ,MRG11 ,MRG12 ,ICEFLERR ,ICENOECC ;
  wire  DCER ,DSER ,DWWR ,DWED ,DMRG00 ,DMRG01 ,DMRG10 ,DMRG11 ;
  wire  DMRG12 ,DREAD ,AF19 ,AF18 ,AF13 ,AF12 ,AF11 ,AF10 ;
  wire  AF1 ,AF0 ,OCDMOD ,CLK60MHZ ,CLK30MHZ_GB ,GDRAMWR ,PSEUDOON10 ,PERISVIB ;
  wire  PSEUDOON1 ,SVMODI ,SVMODIPERI1 ,SVMODIPERI2 ,STBRELESV ,PONRESB ,CPUPRCLK3 ,CPURCLK3 ;
  wire  CPUTMCLK ,CPUMCLK ,CPUTSCLK ,CPUSCLK ,POCRESB ,VDDLEV0 ,VDDLEV1 ,VDDLEV2 ;
  wire  VDDLEV3 ,VDDLEV4 ,VDDLEV5 ,VDDLEV6 ,VDDLEV7 ,USBIFWR ,PSEUDOON0 ,PSEUDOON8 ;
  wire  RESFB5V ,ICEWR ,ICEIFA0 ,ICEIFA1 ,ICEIFA5 ,ICEIFA6 ,ICEIFA7 ,ICEIFA8 ;
  wire  ICEIFA9 ,ICEIFA10 ,ICEIFA11 ,ICEIFA12 ,ICEIFA20 ,ICEIFA13 ,ICEIFA21 ,ICEIFA14 ;
  wire  ICEIFA22 ,ICEIFA30 ,ICEIFA15 ,ICEIFA23 ,ICEIFA31 ,ICEIFA16 ,ICEIFA24 ,ICEIFA17 ;
  wire  ICEIFA25 ,ICEIFA18 ,ICEIFA26 ,ICEIFA19 ,ICEIFA27 ,ICEIFA28 ,ICEIFA29 ,ICEDI0 ;
  wire  ICEDI1 ,ICEDI10 ,ICEDI11 ,ICEDI12 ,ICEDI20 ,ICEDI13 ,ICEDI21 ,ICEDOP0 ;
  wire  ICEDOP1 ,ICEDOP2 ,ICEDOP3 ,ICEDOP4 ,ICEDOP5 ,ICEDOP6 ,ICEDOP7 ,ICEDOP8 ;
  wire  ICEDOP9 ,ICEDOP10 ,ICEDOP11 ,ICEDOP12 ,ICEDOP20 ,ICEDOP13 ,ICEDOP21 ,ICEDOP14 ;
  wire  ICEDOP22 ,ICEDOP30 ,ICEDOP15 ,ICEDOP23 ,ICEDOP31 ,ICEDOP16 ,ICEDOP24 ,ICEDOP17 ;
  wire  ICEDOP25 ,ICEDOP18 ,ICEDOP26 ,ICEDOP19 ,ICEDOP27 ,ICEDOP28 ,ICEDOP29 ,STOPZ ;
  wire  P00ENO ,P01ENO ,P02ENO ,P10ENO ,P03ENO ,P11ENO ,P04ENO ,P12ENO ;
  wire  P20ENO ,P05ENO ,P13ENO ,P21ENO ,P06ENO ,P14ENO ,P22ENO ,P30ENO ;
  wire  P00DOUT ,P01DOUT ,P02DOUT ,P10DOUT ,P03DOUT ,P11DOUT ,P04DOUT ,P12DOUT ;
  wire  P20DOUT ,ADDRTD2 ,P05DOUT ,P13DOUT ,P21DOUT ,P06DOUT ,P14DOUT ,P22DOUT ;
  wire  P30DOUT ,P00ENI ,P01ENI ,P02ENI ,P10ENI ,P03ENI ,P11ENI ,P04ENI ;
  wire  P12ENI ,P20ENI ,P05ENI ,P13ENI ,P21ENI ,P06ENI ,P14ENI ,P22ENI ;
  wire  P30ENI ,P00DIN ,P01DIN ,P02DIN ,P10DIN ,P03DIN ,P11DIN ,P04DIN ;
  wire  P12DIN ,P20DIN ,P05DIN ,P13DIN ,P21DIN ,P06DIN ,P14DIN ,P22DIN ;
  wire  P30DIN ,P01SELIN ,P03SELIN ,P11SELIN ,P04SELIN ,P15ENO ,P23ENO ,P31ENO ;
  wire  P16ENO ,P24ENO ,P40ENO ,P17ENO ,P25ENO ,P41ENO ,P15DOUT ,P23DOUT ;
  wire  P31DOUT ,P16DOUT ,P24DOUT ,P40DOUT ,P17DOUT ,P25DOUT ,P41DOUT ,P15ENI ;
  wire  P23ENI ,P31ENI ,P16ENI ,P24ENI ,P40ENI ,P17ENI ,P25ENI ,P41ENI ;
  wire  P15DIN ,P23DIN ,P31DIN ,P16DIN ,P24DIN ,P40DIN ,P17DIN ,P25DIN ;
  wire  P41DIN ,P10SELIN ,P13SELIN ,P14SELIN ,P15SELIN ,P16SELIN ,P17SELIN ,P26ENO ;
  wire  P42ENO ,P50ENO ,P27ENO ,P43ENO ,P51ENO ,P26DOUT ,P42DOUT ,P50DOUT ;
  wire  P27DOUT ,P43DOUT ,P51DOUT ,P26ENI ,P42ENI ,P50ENI ,P27ENI ,P43ENI ;
  wire  P51ENI ,P26DIN ,P42DIN ,P50DIN ,P27DIN ,P43DIN ,P51DIN ,P52ENO ;
  wire  P60ENO ,P53ENO ,P61ENO ,DGEN07 ,P54ENO ,P62ENO ,P70ENO ,P55ENO ;
  wire  P63ENO ,P71ENO ,P52DOUT ,P60DOUT ,P53DOUT ,P61DOUT ,P54DOUT ,P62DOUT ;
  wire  P70DOUT ,P55DOUT ,P63DOUT ,P71DOUT ,P52ENI ,P60ENI ,P53ENI ,P61ENI ;
  wire  DGEN01 ,P54ENI ,P62ENI ,P70ENI ,P55ENI ,P63ENI ,P71ENI ,P52DIN ;
  wire  P60DIN ,P53DIN ,P61DIN ,P54DIN ,P62DIN ,P70DIN ,DGEN00 ,P55DIN ;
  wire  P63DIN ,P71DIN ,P55SELIN ,P72ENO ,P73ENO ,P74ENO ,P75ENO ,P77ENO ;
  wire  P72DOUT ,P73DOUT ,P74DOUT ,P75DOUT ,P76DOUT ,P77DOUT ,P72ENI ,P73ENI ;
  wire  P74ENI ,P75ENI ,P76ENI ,P72DIN ,P73DIN ,P75DIN ,P76DIN ,P120ENO ;
  wire  P120DOUT ,P120ENI ,P120DIN ,P130ENO ,P130DOUT ,P137ENI ,P137DIN ,P140ENO ;
  wire  P141ENO ,P146ENO ,P147ENO ,P140DOUT ,P141DOUT ,P146DOUT ,P147DOUT ,P140ENI ;
  wire  P141ENI ,P146ENI ,P147ENI ,P140DIN ,P141DIN ,P146DIN ,P147DIN ,P00PUON ;
  wire  P01PUON ,P02PUON ,P10PUON ,P03PUON ,P11PUON ,P04PUON ,P12PUON ,P06PUON ;
  wire  P14PUON ,P30PUON ,P15PUON ,P31PUON ,P16PUON ,P40PUON ,P17PUON ,P41PUON ;
  wire  P43PUON ,P51PUON ,P52PUON ,P53PUON ,P54PUON ,P70PUON ,P55PUON ,P71PUON ;
  wire  P72PUON ,P75PUON ,P76PUON ,P77PUON ,P120PUON ,P140PUON ,P141PUON ,P146PUON ;
  wire  P147PUON ,PIO137 ,PSEUDOANI09 ,PSEUDOANI17 ,PSEUDOANI08 ,PSEUDOANI16 ,PSEUDOANI07 ,PSEUDOANI15 ;
  wire  PSEUDOANI06 ,PSEUDOANI14 ,PSEUDOANI05 ,PSEUDOANI13 ,PSEUDOANI04 ,PSEUDOANI12 ,PSEUDOANI03 ,PSEUDOANI11 ;
  wire  PSEUDOANI02 ,PSEUDOANI10 ,PSEUDOANI01 ,PSEUDOANI00 ,PSEUDOANI19 ,PSEUDOANI18 ,ADVSELMOD0_I ,ADVSELMOD1_I ;
  wire  DGEN06 ,DGEN05 ,DGEN04 ,DGEN03 ,DGEN02 ,CLK60MHZLOCK ,CPURCLK1 ,CPURCLK2 ;
  wire  SVMODOPBRK ,PSEUDOON31 ,PSEUDOON23 ,PSEUDOON15 ,PSEUDOON30 ,PSEUDOON22 ,PSEUDOON14 ,PSEUDOON29 ;
  wire  PSEUDOON28 ,PSEUDOON27 ,PSEUDOON19 ,PSEUDOON26 ,PSEUDOON18 ,PSEUDOON25 ,PSEUDOON17 ,PSEUDOON24 ;
  wire  PSEUDOON16 ,PSEUDOON21 ,PSEUDOON13 ,PSEUDOON20 ,PSEUDOON12 ,PSEUDOON11 ,PSEUDOON9 ,ICEMSKWAIT ;
  wire  ICEMSKTRAP ,ICEMSKRETRY ,IDVER31 ,IDVER23 ,IDVER15 ,IDVER30 ,IDVER22 ,IDVER14 ;
  wire  IDVER29 ,IDVER28 ,IDVER27 ,IDVER19 ,IDVER26 ,IDVER18 ,IDVER25 ,IDVER17 ;
  wire  IDVER24 ,IDVER16 ,IDVER21 ,IDVER13 ,IDVER20 ,IDVER12 ,IDVER11 ,IDVER10 ;
  wire  IDVER9 ,IDVER8 ,IDVER7 ,IDVER6 ,IDVER5 ,IDVER4 ,IDVER3 ,IDVER2 ;
  wire  IDVER1 ,IDVER0 ,ADDRTD144 ,ADDRTD136 ,ADDRTD128 ,ADDRTD143 ,ADDRTD135 ,ADDRTD127 ;
  wire  ADDRTD119 ,ADDRTD142 ,ADDRTD134 ,ADDRTD126 ,ADDRTD118 ,ADDRTD141 ,ADDRTD133 ,ADDRTD125 ;
  wire  ADDRTD117 ,ADDRTD109 ,ADDRTD140 ,ADDRTD132 ,ADDRTD124 ,ADDRTD116 ,ADDRTD108 ,ADDRTD139 ;
  wire  ADDRTD138 ,ADDRTD137 ,ADDRTD129 ,ADDRTD131 ,ADDRTD123 ,ADDRTD115 ,ADDRTD107 ,ADDRTD130 ;
  wire  ADDRTD122 ,ADDRTD114 ,ADDRTD106 ,ADDRTD121 ,ADDRTD113 ,ADDRTD105 ,ADDRTD120 ,ADDRTD112 ;
  wire  ADDRTD104 ,ADDRTD111 ,ADDRTD103 ,ADDRTD110 ,ADDRTD102 ,ADDRTD101 ,ADDRTD100 ,ADDRTD99 ;
  wire  ADDRTD98 ,ADDRTD97 ,ADDRTD89 ,ADDRTD96 ,ADDRTD88 ,ADDRTD95 ,ADDRTD87 ,ADDRTD79 ;
  wire  ADDRTD94 ,ADDRTD86 ,ADDRTD78 ,ADDRTD93 ,ADDRTD85 ,ADDRTD77 ,ADDRTD69 ,ADDRTD92 ;
  wire  ADDRTD84 ,ADDRTD76 ,ADDRTD68 ,ADDRTD91 ,ADDRTD83 ,ADDRTD75 ,ADDRTD67 ,ADDRTD59 ;
  wire  ADDRTD90 ,ADDRTD82 ,ADDRTD74 ,ADDRTD66 ,ADDRTD58 ,ADDRTD81 ,ADDRTD73 ,ADDRTD65 ;
  wire  ADDRTD57 ,ADDRTD49 ,ADDRTD80 ,ADDRTD72 ,ADDRTD64 ,ADDRTD56 ,ADDRTD48 ,ADDRTD71 ;
  wire  ADDRTD63 ,ADDRTD55 ,ADDRTD47 ,ADDRTD39 ,ADDRTD70 ,ADDRTD62 ,ADDRTD54 ,ADDRTD46 ;
  wire  ADDRTD38 ,ADDRTD61 ,ADDRTD53 ,ADDRTD45 ,ADDRTD37 ,ADDRTD29 ,ADDRTD60 ,ADDRTD52 ;
  wire  ADDRTD44 ,ADDRTD36 ,ADDRTD28 ,ADDRTD51 ,ADDRTD43 ,ADDRTD35 ,ADDRTD27 ,ADDRTD19 ;
  wire  ADDRTD50 ,ADDRTD42 ,ADDRTD34 ,ADDRTD26 ,ADDRTD18 ,ADDRTD41 ,ADDRTD33 ,ADDRTD25 ;
  wire  ADDRTD17 ,ADDRTD40 ,ADDRTD32 ,ADDRTD24 ,ADDRTD16 ,ADDRTD31 ,ADDRTD23 ,ADDRTD15 ;
  wire  ADDRTD30 ,ADDRTD22 ,ADDRTD14 ,ADDRTD21 ,ADDRTD13 ,ADDRTD20 ,ADDRTD12 ,ADDRTD11 ;
  wire  ADDRTD10 ,ADDRTD9 ,ADDRTD8 ,ADDRTD7 ,ADDRTD6 ,ADDRTD5 ,ADDRTD4 ,ADDRTD3 ;
  wire  ADDRTD1 ,ADDRPINRD ,ADDRPINMD ,ADDRPINLV ,DDIS_OUT ,DRDCLKP1_OUT ,DWWR_OUT ,DCER_OUT ;
  wire  DSER_OUT ,DMRG00_OUT ,DMRG01_OUT ,DMRG10_OUT ,DMRG11_OUT ,DMRG12_OUT ,DREAD_OUT ,DFCLK_OUT ;

  TBCLL pulldown0 ( pull_down0 ) ;
  TBCLL pulldown1 ( pull_down1 ) ;
  TBCLL pulldown2 ( pull_down2 ) ;
  TBCLL pulldown3 ( pull_down3 ) ;
  TBCLL pulldown4 ( pull_down4 ) ;
  TBCLL pulldown5 ( pull_down5 ) ;
  TBCLL pulldown6 ( pull_down6 ) ;
  TBCLL pulldown7 ( pull_down7 ) ;
  TBCLL pulldown8 ( pull_down8 ) ;
  TBCLL pulldown9 ( pull_down9 ) ;
  TBCLL pulldown10 ( pull_down10 ) ;
  TBCLL pulldown11 ( pull_down11 ) ;
  TBCLL pulldown12 ( pull_down12 ) ;
  TBCLL pulldown20 ( pull_down20 ) ;
  TBCLL pulldown13 ( pull_down13 ) ;
  TBCLL pulldown21 ( pull_down21 ) ;
  TBCLL pulldown14 ( pull_down14 ) ;
  TBCLL pulldown22 ( pull_down22 ) ;
  TBCLL pulldown30 ( pull_down30 ) ;
  TBCLL pulldown15 ( pull_down15 ) ;
  TBCLL pulldown23 ( pull_down23 ) ;
  TBCLL pulldown31 ( pull_down31 ) ;
  TBCLL pulldown16 ( pull_down16 ) ;
  TBCLL pulldown24 ( pull_down24 ) ;
  TBCLL pulldown32 ( pull_down32 ) ;
  TBCLL pulldown40 ( pull_down40 ) ;
  TBCLL pulldown17 ( pull_down17 ) ;
  TBCLL pulldown25 ( pull_down25 ) ;
  TBCLL pulldown33 ( pull_down33 ) ;
  TBCLL pulldown41 ( pull_down41 ) ;
  TBCLL pulldown18 ( pull_down18 ) ;
  TBCLL pulldown26 ( pull_down26 ) ;
  TBCLL pulldown34 ( pull_down34 ) ;
  TBCLL pulldown42 ( pull_down42 ) ;
  TBCLL pulldown50 ( pull_down50 ) ;
  TBCLL pulldown19 ( pull_down19 ) ;
  TBCLL pulldown27 ( pull_down27 ) ;
  TBCLL pulldown35 ( pull_down35 ) ;
  TBCLL pulldown43 ( pull_down43 ) ;
  TBCLL pulldown51 ( pull_down51 ) ;
  TBCLL pulldown28 ( pull_down28 ) ;
  TBCLL pulldown36 ( pull_down36 ) ;
  TBCLL pulldown44 ( pull_down44 ) ;
  TBCLL pulldown52 ( pull_down52 ) ;
  TBCLL pulldown60 ( pull_down60 ) ;
  TBCLL pulldown29 ( pull_down29 ) ;
  TBCLL pulldown37 ( pull_down37 ) ;
  TBCLL pulldown45 ( pull_down45 ) ;
  TBCLL pulldown53 ( pull_down53 ) ;
  TBCLL pulldown61 ( pull_down61 ) ;
  TBCLL pulldown38 ( pull_down38 ) ;
  TBCLL pulldown46 ( pull_down46 ) ;
  TBCLL pulldown54 ( pull_down54 ) ;
  TBCLL pulldown62 ( pull_down62 ) ;
  TBCLL pulldown70 ( pull_down70 ) ;
  TBCLL pulldown39 ( pull_down39 ) ;
  TBCLL pulldown47 ( pull_down47 ) ;
  TBCLL pulldown55 ( pull_down55 ) ;
  TBCLL pulldown63 ( pull_down63 ) ;
  TBCLL pulldown71 ( pull_down71 ) ;
  TBCLL pulldown48 ( pull_down48 ) ;
  TBCLL pulldown56 ( pull_down56 ) ;
  TBCLL pulldown64 ( pull_down64 ) ;
  TBCLL pulldown72 ( pull_down72 ) ;
  TBCLL pulldown80 ( pull_down80 ) ;
  TBCLL pulldown49 ( pull_down49 ) ;
  TBCLL pulldown57 ( pull_down57 ) ;
  TBCLL pulldown65 ( pull_down65 ) ;
  TBCLL pulldown73 ( pull_down73 ) ;
  TBCLL pulldown81 ( pull_down81 ) ;
  TBCLL pulldown58 ( pull_down58 ) ;
  TBCLL pulldown66 ( pull_down66 ) ;
  TBCLL pulldown74 ( pull_down74 ) ;
  TBCLL pulldown82 ( pull_down82 ) ;
  TBCLL pulldown90 ( pull_down90 ) ;
  TBCLL pulldown59 ( pull_down59 ) ;
  TBCLL pulldown67 ( pull_down67 ) ;
  TBCLL pulldown75 ( pull_down75 ) ;
  TBCLL pulldown83 ( pull_down83 ) ;
  TBCLL pulldown91 ( pull_down91 ) ;
  TBCLL pulldown68 ( pull_down68 ) ;
  TBCLL pulldown76 ( pull_down76 ) ;
  TBCLL pulldown84 ( pull_down84 ) ;
  TBCLL pulldown92 ( pull_down92 ) ;
  TBCLL pulldown69 ( pull_down69 ) ;
  TBCLL pulldown77 ( pull_down77 ) ;
  TBCLL pulldown85 ( pull_down85 ) ;
  TBCLL pulldown93 ( pull_down93 ) ;
  TBCLL pulldown78 ( pull_down78 ) ;
  TBCLL pulldown86 ( pull_down86 ) ;
  TBCLL pulldown94 ( pull_down94 ) ;
  TBCLL pulldown79 ( pull_down79 ) ;
  TBCLL pulldown87 ( pull_down87 ) ;
  TBCLL pulldown95 ( pull_down95 ) ;
  TBCLL pulldown88 ( pull_down88 ) ;
  TBCLL pulldown96 ( pull_down96 ) ;
  TBCLL pulldown89 ( pull_down89 ) ;
  TBCLL pulldown97 ( pull_down97 ) ;
  TBCLL pulldown98 ( pull_down98 ) ;
  TBCLL pulldown99 ( pull_down99 ) ;
  TBCLL pulldown100 ( pull_down100 ) ;
  TBCLL pulldown101 ( pull_down101 ) ;
  TBCLL pulldown102 ( pull_down102 ) ;
  TBCLL pulldown110 ( pull_down110 ) ;
  TBCLL pulldown103 ( pull_down103 ) ;
  TBCLL pulldown111 ( pull_down111 ) ;
  TBCLL pulldown104 ( pull_down104 ) ;
  TBCLL pulldown112 ( pull_down112 ) ;
  TBCLL pulldown120 ( pull_down120 ) ;
  TBCLL pulldown200 ( pull_down200 ) ;
  TBCLL pulldown105 ( pull_down105 ) ;
  TBCLL pulldown113 ( pull_down113 ) ;
  TBCLL pulldown121 ( pull_down121 ) ;
  TBCLL pulldown201 ( pull_down201 ) ;
  TBCLL pulldown106 ( pull_down106 ) ;
  TBCLL pulldown114 ( pull_down114 ) ;
  TBCLL pulldown122 ( pull_down122 ) ;
  TBCLL pulldown130 ( pull_down130 ) ;
  TBCLL pulldown202 ( pull_down202 ) ;
  TBCLL pulldown210 ( pull_down210 ) ;
  TBCLL pulldown107 ( pull_down107 ) ;
  TBCLL pulldown115 ( pull_down115 ) ;
  TBCLL pulldown123 ( pull_down123 ) ;
  TBCLL pulldown131 ( pull_down131 ) ;
  TBCLL pulldown203 ( pull_down203 ) ;
  TBCLL pulldown211 ( pull_down211 ) ;
  TBCLL pulldown108 ( pull_down108 ) ;
  TBCLL pulldown116 ( pull_down116 ) ;
  TBCLL pulldown124 ( pull_down124 ) ;
  TBCLL pulldown132 ( pull_down132 ) ;
  TBCLL pulldown140 ( pull_down140 ) ;
  TBCLL pulldown204 ( pull_down204 ) ;
  TBCLL pulldown212 ( pull_down212 ) ;
  TBCLL pulldown220 ( pull_down220 ) ;
  TBCLL pulldown300 ( pull_down300 ) ;
  TBCLL pulldown109 ( pull_down109 ) ;
  TBCLL pulldown117 ( pull_down117 ) ;
  TBCLL pulldown125 ( pull_down125 ) ;
  TBCLL pulldown133 ( pull_down133 ) ;
  TBCLL pulldown141 ( pull_down141 ) ;
  TBCLL pulldown205 ( pull_down205 ) ;
  TBCLL pulldown213 ( pull_down213 ) ;
  TBCLL pulldown221 ( pull_down221 ) ;
  TBCLL pulldown301 ( pull_down301 ) ;
  TBCLL pulldown118 ( pull_down118 ) ;
  TBCLL pulldown126 ( pull_down126 ) ;
  TBCLL pulldown134 ( pull_down134 ) ;
  TBCLL pulldown142 ( pull_down142 ) ;
  TBCLL pulldown150 ( pull_down150 ) ;
  TBCLL pulldown206 ( pull_down206 ) ;
  TBCLL pulldown214 ( pull_down214 ) ;
  TBCLL pulldown222 ( pull_down222 ) ;
  TBCLL pulldown230 ( pull_down230 ) ;
  TBCLL pulldown302 ( pull_down302 ) ;
  TBCLL pulldown310 ( pull_down310 ) ;
  TBCLL pulldown119 ( pull_down119 ) ;
  TBCLL pulldown127 ( pull_down127 ) ;
  TBCLL pulldown135 ( pull_down135 ) ;
  TBCLL pulldown143 ( pull_down143 ) ;
  TBCLL pulldown151 ( pull_down151 ) ;
  TBCLL pulldown207 ( pull_down207 ) ;
  TBCLL pulldown215 ( pull_down215 ) ;
  TBCLL pulldown223 ( pull_down223 ) ;
  TBCLL pulldown231 ( pull_down231 ) ;
  TBCLL pulldown303 ( pull_down303 ) ;
  TBCLL pulldown311 ( pull_down311 ) ;
  TBCLL pulldown128 ( pull_down128 ) ;
  TBCLL pulldown136 ( pull_down136 ) ;
  TBCLL pulldown144 ( pull_down144 ) ;
  TBCLL pulldown152 ( pull_down152 ) ;
  TBCLL pulldown160 ( pull_down160 ) ;
  TBCLL pulldown208 ( pull_down208 ) ;
  TBCLL pulldown216 ( pull_down216 ) ;
  TBCLL pulldown224 ( pull_down224 ) ;
  TBCLL pulldown232 ( pull_down232 ) ;
  TBCLL pulldown240 ( pull_down240 ) ;
  TBCLL pulldown304 ( pull_down304 ) ;
  TBCLL pulldown312 ( pull_down312 ) ;
  TBCLL pulldown320 ( pull_down320 ) ;
  TBCLL pulldown400 ( pull_down400 ) ;
  TBCLL pulldown129 ( pull_down129 ) ;
  TBCLL pulldown137 ( pull_down137 ) ;
  TBCLL pulldown145 ( pull_down145 ) ;
  TBCLL pulldown153 ( pull_down153 ) ;
  TBCLL pulldown161 ( pull_down161 ) ;
  TBCLL pulldown209 ( pull_down209 ) ;
  TBCLL pulldown217 ( pull_down217 ) ;
  TBCLL pulldown225 ( pull_down225 ) ;
  TBCLL pulldown233 ( pull_down233 ) ;
  TBCLL pulldown241 ( pull_down241 ) ;
  TBCLL pulldown305 ( pull_down305 ) ;
  TBCLL pulldown313 ( pull_down313 ) ;
  TBCLL pulldown321 ( pull_down321 ) ;
  TBCLL pulldown401 ( pull_down401 ) ;
  TBCLL pulldown138 ( pull_down138 ) ;
  TBCLL pulldown146 ( pull_down146 ) ;
  TBCLL pulldown154 ( pull_down154 ) ;
  TBCLL pulldown162 ( pull_down162 ) ;
  TBCLL pulldown170 ( pull_down170 ) ;
  TBCLL pulldown218 ( pull_down218 ) ;
  TBCLL pulldown226 ( pull_down226 ) ;
  TBCLL pulldown234 ( pull_down234 ) ;
  TBCLL pulldown242 ( pull_down242 ) ;
  TBCLL pulldown250 ( pull_down250 ) ;
  TBCLL pulldown306 ( pull_down306 ) ;
  TBCLL pulldown314 ( pull_down314 ) ;
  TBCLL pulldown322 ( pull_down322 ) ;
  TBCLL pulldown330 ( pull_down330 ) ;
  TBCLL pulldown402 ( pull_down402 ) ;
  TBCLL pulldown410 ( pull_down410 ) ;
  TBCLL pulldown139 ( pull_down139 ) ;
  TBCLL pulldown147 ( pull_down147 ) ;
  TBCLL pulldown155 ( pull_down155 ) ;
  TBCLL pulldown163 ( pull_down163 ) ;
  TBCLL pulldown171 ( pull_down171 ) ;
  TBCLL pulldown219 ( pull_down219 ) ;
  TBCLL pulldown227 ( pull_down227 ) ;
  TBCLL pulldown235 ( pull_down235 ) ;
  TBCLL pulldown243 ( pull_down243 ) ;
  TBCLL pulldown251 ( pull_down251 ) ;
  TBCLL pulldown307 ( pull_down307 ) ;
  TBCLL pulldown315 ( pull_down315 ) ;
  TBCLL pulldown323 ( pull_down323 ) ;
  TBCLL pulldown331 ( pull_down331 ) ;
  TBCLL pulldown403 ( pull_down403 ) ;
  TBCLL pulldown411 ( pull_down411 ) ;
  TBCLL pulldown148 ( pull_down148 ) ;
  TBCLL pulldown156 ( pull_down156 ) ;
  TBCLL pulldown164 ( pull_down164 ) ;
  TBCLL pulldown172 ( pull_down172 ) ;
  TBCLL pulldown180 ( pull_down180 ) ;
  TBCLL pulldown228 ( pull_down228 ) ;
  TBCLL pulldown236 ( pull_down236 ) ;
  TBCLL pulldown244 ( pull_down244 ) ;
  TBCLL pulldown252 ( pull_down252 ) ;
  TBCLL pulldown260 ( pull_down260 ) ;
  TBCLL pulldown308 ( pull_down308 ) ;
  TBCLL pulldown316 ( pull_down316 ) ;
  TBCLL pulldown324 ( pull_down324 ) ;
  TBCLL pulldown332 ( pull_down332 ) ;
  TBCLL pulldown340 ( pull_down340 ) ;
  TBCLL pulldown404 ( pull_down404 ) ;
  TBCLL pulldown412 ( pull_down412 ) ;
  TBCLL pulldown420 ( pull_down420 ) ;
  TBCLL pulldown500 ( pull_down500 ) ;
  TBCLL pulldown149 ( pull_down149 ) ;
  TBCLL pulldown157 ( pull_down157 ) ;
  TBCLL pulldown165 ( pull_down165 ) ;
  TBCLL pulldown173 ( pull_down173 ) ;
  TBCLL pulldown181 ( pull_down181 ) ;
  TBCLL pulldown229 ( pull_down229 ) ;
  TBCLL pulldown237 ( pull_down237 ) ;
  TBCLL pulldown245 ( pull_down245 ) ;
  TBCLL pulldown253 ( pull_down253 ) ;
  TBCLL pulldown261 ( pull_down261 ) ;
  TBCLL pulldown309 ( pull_down309 ) ;
  TBCLL pulldown317 ( pull_down317 ) ;
  TBCLL pulldown325 ( pull_down325 ) ;
  TBCLL pulldown333 ( pull_down333 ) ;
  TBCLL pulldown341 ( pull_down341 ) ;
  TBCLL pulldown405 ( pull_down405 ) ;
  TBCLL pulldown413 ( pull_down413 ) ;
  TBCLL pulldown421 ( pull_down421 ) ;
  TBCLL pulldown501 ( pull_down501 ) ;
  TBCLL pulldown158 ( pull_down158 ) ;
  TBCLL pulldown166 ( pull_down166 ) ;
  TBCLL pulldown174 ( pull_down174 ) ;
  TBCLL pulldown182 ( pull_down182 ) ;
  TBCLL pulldown190 ( pull_down190 ) ;
  TBCLL pulldown238 ( pull_down238 ) ;
  TBCLL pulldown246 ( pull_down246 ) ;
  TBCLL pulldown254 ( pull_down254 ) ;
  TBCLL pulldown262 ( pull_down262 ) ;
  TBCLL pulldown270 ( pull_down270 ) ;
  TBCLL pulldown318 ( pull_down318 ) ;
  TBCLL pulldown326 ( pull_down326 ) ;
  TBCLL pulldown334 ( pull_down334 ) ;
  TBCLL pulldown342 ( pull_down342 ) ;
  TBCLL pulldown350 ( pull_down350 ) ;
  TBCLL pulldown406 ( pull_down406 ) ;
  TBCLL pulldown414 ( pull_down414 ) ;
  TBCLL pulldown422 ( pull_down422 ) ;
  TBCLL pulldown430 ( pull_down430 ) ;
  TBCLL pulldown502 ( pull_down502 ) ;
  TBCLL pulldown510 ( pull_down510 ) ;
  TBCLL pulldown159 ( pull_down159 ) ;
  TBCLL pulldown167 ( pull_down167 ) ;
  TBCLL pulldown175 ( pull_down175 ) ;
  TBCLL pulldown183 ( pull_down183 ) ;
  TBCLL pulldown191 ( pull_down191 ) ;
  TBCLL pulldown239 ( pull_down239 ) ;
  TBCLL pulldown247 ( pull_down247 ) ;
  TBCLL pulldown255 ( pull_down255 ) ;
  TBCLL pulldown263 ( pull_down263 ) ;
  TBCLL pulldown271 ( pull_down271 ) ;
  TBCLL pulldown319 ( pull_down319 ) ;
  TBCLL pulldown327 ( pull_down327 ) ;
  TBCLL pulldown335 ( pull_down335 ) ;
  TBCLL pulldown343 ( pull_down343 ) ;
  TBCLL pulldown351 ( pull_down351 ) ;
  TBCLL pulldown407 ( pull_down407 ) ;
  TBCLL pulldown415 ( pull_down415 ) ;
  TBCLL pulldown423 ( pull_down423 ) ;
  TBCLL pulldown431 ( pull_down431 ) ;
  TBCLL pulldown503 ( pull_down503 ) ;
  TBCLL pulldown511 ( pull_down511 ) ;
  TBCLL pulldown168 ( pull_down168 ) ;
  TBCLL pulldown176 ( pull_down176 ) ;
  TBCLL pulldown184 ( pull_down184 ) ;
  TBCLL pulldown192 ( pull_down192 ) ;
  TBCLL pulldown248 ( pull_down248 ) ;
  TBCLL pulldown256 ( pull_down256 ) ;
  TBCLL pulldown264 ( pull_down264 ) ;
  TBCLL pulldown272 ( pull_down272 ) ;
  TBCLL pulldown280 ( pull_down280 ) ;
  TBCLL pulldown328 ( pull_down328 ) ;
  TBCLL pulldown336 ( pull_down336 ) ;
  TBCLL pulldown344 ( pull_down344 ) ;
  TBCLL pulldown352 ( pull_down352 ) ;
  TBCLL pulldown360 ( pull_down360 ) ;
  TBCLL pulldown408 ( pull_down408 ) ;
  TBCLL pulldown416 ( pull_down416 ) ;
  TBCLL pulldown424 ( pull_down424 ) ;
  TBCLL pulldown432 ( pull_down432 ) ;
  TBCLL pulldown440 ( pull_down440 ) ;
  TBCLL pulldown504 ( pull_down504 ) ;
  TBCLL pulldown512 ( pull_down512 ) ;
  TBCLL pulldown520 ( pull_down520 ) ;
  TBCLL pulldown600 ( pull_down600 ) ;
  TBCLL pulldown169 ( pull_down169 ) ;
  TBCLL pulldown177 ( pull_down177 ) ;
  TBCLL pulldown185 ( pull_down185 ) ;
  TBCLL pulldown193 ( pull_down193 ) ;
  TBCLL pulldown249 ( pull_down249 ) ;
  TBCLL pulldown257 ( pull_down257 ) ;
  TBCLL pulldown265 ( pull_down265 ) ;
  TBCLL pulldown273 ( pull_down273 ) ;
  TBCLL pulldown281 ( pull_down281 ) ;
  TBCLL pulldown329 ( pull_down329 ) ;
  TBCLL pulldown337 ( pull_down337 ) ;
  TBCLL pulldown345 ( pull_down345 ) ;
  TBCLL pulldown353 ( pull_down353 ) ;
  TBCLL pulldown361 ( pull_down361 ) ;
  TBCLL pulldown409 ( pull_down409 ) ;
  TBCLL pulldown417 ( pull_down417 ) ;
  TBCLL pulldown425 ( pull_down425 ) ;
  TBCLL pulldown433 ( pull_down433 ) ;
  TBCLL pulldown441 ( pull_down441 ) ;
  TBCLL pulldown505 ( pull_down505 ) ;
  TBCLL pulldown513 ( pull_down513 ) ;
  TBCLL pulldown521 ( pull_down521 ) ;
  TBCLL pulldown601 ( pull_down601 ) ;
  TBCLL pulldown178 ( pull_down178 ) ;
  TBCLL pulldown186 ( pull_down186 ) ;
  TBCLL pulldown194 ( pull_down194 ) ;
  TBCLL pulldown258 ( pull_down258 ) ;
  TBCLL pulldown266 ( pull_down266 ) ;
  TBCLL pulldown274 ( pull_down274 ) ;
  TBCLL pulldown282 ( pull_down282 ) ;
  TBCLL pulldown290 ( pull_down290 ) ;
  TBCLL pulldown338 ( pull_down338 ) ;
  TBCLL pulldown346 ( pull_down346 ) ;
  TBCLL pulldown354 ( pull_down354 ) ;
  TBCLL pulldown362 ( pull_down362 ) ;
  TBCLL pulldown370 ( pull_down370 ) ;
  TBCLL pulldown418 ( pull_down418 ) ;
  TBCLL pulldown426 ( pull_down426 ) ;
  TBCLL pulldown434 ( pull_down434 ) ;
  TBCLL pulldown442 ( pull_down442 ) ;
  TBCLL pulldown450 ( pull_down450 ) ;
  TBCLL pulldown506 ( pull_down506 ) ;
  TBCLL pulldown514 ( pull_down514 ) ;
  TBCLL pulldown522 ( pull_down522 ) ;
  TBCLL pulldown530 ( pull_down530 ) ;
  TBCLL pulldown602 ( pull_down602 ) ;
  TBCLL pulldown610 ( pull_down610 ) ;
  TBCLL pulldown179 ( pull_down179 ) ;
  TBCLL pulldown187 ( pull_down187 ) ;
  TBCLL pulldown195 ( pull_down195 ) ;
  TBCLL pulldown259 ( pull_down259 ) ;
  TBCLL pulldown267 ( pull_down267 ) ;
  TBCLL pulldown275 ( pull_down275 ) ;
  TBCLL pulldown283 ( pull_down283 ) ;
  TBCLL pulldown291 ( pull_down291 ) ;
  TBCLL pulldown339 ( pull_down339 ) ;
  TBCLL pulldown347 ( pull_down347 ) ;
  TBCLL pulldown355 ( pull_down355 ) ;
  TBCLL pulldown363 ( pull_down363 ) ;
  TBCLL pulldown371 ( pull_down371 ) ;
  TBCLL pulldown419 ( pull_down419 ) ;
  TBCLL pulldown427 ( pull_down427 ) ;
  TBCLL pulldown435 ( pull_down435 ) ;
  TBCLL pulldown443 ( pull_down443 ) ;
  TBCLL pulldown451 ( pull_down451 ) ;
  TBCLL pulldown507 ( pull_down507 ) ;
  TBCLL pulldown515 ( pull_down515 ) ;
  TBCLL pulldown523 ( pull_down523 ) ;
  TBCLL pulldown531 ( pull_down531 ) ;
  TBCLL pulldown603 ( pull_down603 ) ;
  TBCLL pulldown611 ( pull_down611 ) ;
  TBCLL pulldown188 ( pull_down188 ) ;
  TBCLL pulldown196 ( pull_down196 ) ;
  TBCLL pulldown268 ( pull_down268 ) ;
  TBCLL pulldown276 ( pull_down276 ) ;
  TBCLL pulldown284 ( pull_down284 ) ;
  TBCLL pulldown292 ( pull_down292 ) ;
  TBCLL pulldown348 ( pull_down348 ) ;
  TBCLL pulldown356 ( pull_down356 ) ;
  TBCLL pulldown364 ( pull_down364 ) ;
  TBCLL pulldown372 ( pull_down372 ) ;
  TBCLL pulldown380 ( pull_down380 ) ;
  TBCLL pulldown428 ( pull_down428 ) ;
  TBCLL pulldown436 ( pull_down436 ) ;
  TBCLL pulldown444 ( pull_down444 ) ;
  TBCLL pulldown452 ( pull_down452 ) ;
  TBCLL pulldown460 ( pull_down460 ) ;
  TBCLL pulldown508 ( pull_down508 ) ;
  TBCLL pulldown516 ( pull_down516 ) ;
  TBCLL pulldown524 ( pull_down524 ) ;
  TBCLL pulldown532 ( pull_down532 ) ;
  TBCLL pulldown540 ( pull_down540 ) ;
  TBCLL pulldown604 ( pull_down604 ) ;
  TBCLL pulldown612 ( pull_down612 ) ;
  TBCLL pulldown620 ( pull_down620 ) ;
  TBCLL pulldown700 ( pull_down700 ) ;
  TBCLL pulldown189 ( pull_down189 ) ;
  TBCLL pulldown197 ( pull_down197 ) ;
  TBCLL pulldown269 ( pull_down269 ) ;
  TBCLL pulldown277 ( pull_down277 ) ;
  TBCLL pulldown285 ( pull_down285 ) ;
  TBCLL pulldown293 ( pull_down293 ) ;
  TBCLL pulldown349 ( pull_down349 ) ;
  TBCLL pulldown357 ( pull_down357 ) ;
  TBCLL pulldown365 ( pull_down365 ) ;
  TBCLL pulldown373 ( pull_down373 ) ;
  TBCLL pulldown381 ( pull_down381 ) ;
  TBCLL pulldown429 ( pull_down429 ) ;
  TBCLL pulldown437 ( pull_down437 ) ;
  TBCLL pulldown445 ( pull_down445 ) ;
  TBCLL pulldown453 ( pull_down453 ) ;
  TBCLL pulldown461 ( pull_down461 ) ;
  TBCLL pulldown509 ( pull_down509 ) ;
  TBCLL pulldown517 ( pull_down517 ) ;
  TBCLL pulldown525 ( pull_down525 ) ;
  TBCLL pulldown533 ( pull_down533 ) ;
  TBCLL pulldown541 ( pull_down541 ) ;
  TBCLL pulldown605 ( pull_down605 ) ;
  TBCLL pulldown613 ( pull_down613 ) ;
  TBCLL pulldown621 ( pull_down621 ) ;
  TBCLL pulldown701 ( pull_down701 ) ;
  TBCLL pulldown198 ( pull_down198 ) ;
  TBCLL pulldown278 ( pull_down278 ) ;
  TBCLL pulldown286 ( pull_down286 ) ;
  TBCLL pulldown294 ( pull_down294 ) ;
  TBCLL pulldown358 ( pull_down358 ) ;
  TBCLL pulldown366 ( pull_down366 ) ;
  TBCLL pulldown374 ( pull_down374 ) ;
  TBCLL pulldown382 ( pull_down382 ) ;
  TBCLL pulldown390 ( pull_down390 ) ;
  TBCLL pulldown438 ( pull_down438 ) ;
  TBCLL pulldown446 ( pull_down446 ) ;
  TBCLL pulldown454 ( pull_down454 ) ;
  TBCLL pulldown462 ( pull_down462 ) ;
  TBCLL pulldown470 ( pull_down470 ) ;
  TBCLL pulldown518 ( pull_down518 ) ;
  TBCLL pulldown526 ( pull_down526 ) ;
  TBCLL pulldown534 ( pull_down534 ) ;
  TBCLL pulldown542 ( pull_down542 ) ;
  TBCLL pulldown550 ( pull_down550 ) ;
  TBCLL pulldown606 ( pull_down606 ) ;
  TBCLL pulldown614 ( pull_down614 ) ;
  TBCLL pulldown622 ( pull_down622 ) ;
  TBCLL pulldown630 ( pull_down630 ) ;
  TBCLL pulldown702 ( pull_down702 ) ;
  TBCLL pulldown710 ( pull_down710 ) ;
  TBCLL pulldown199 ( pull_down199 ) ;
  TBCLL pulldown279 ( pull_down279 ) ;
  TBCLL pulldown287 ( pull_down287 ) ;
  TBCLL pulldown295 ( pull_down295 ) ;
  TBCLL pulldown359 ( pull_down359 ) ;
  TBCLL pulldown367 ( pull_down367 ) ;
  TBCLL pulldown375 ( pull_down375 ) ;
  TBCLL pulldown383 ( pull_down383 ) ;
  TBCLL pulldown391 ( pull_down391 ) ;
  TBCLL pulldown439 ( pull_down439 ) ;
  TBCLL pulldown447 ( pull_down447 ) ;
  TBCLL pulldown455 ( pull_down455 ) ;
  TBCLL pulldown463 ( pull_down463 ) ;
  TBCLL pulldown471 ( pull_down471 ) ;
  TBCLL pulldown519 ( pull_down519 ) ;
  TBCLL pulldown527 ( pull_down527 ) ;
  TBCLL pulldown535 ( pull_down535 ) ;
  TBCLL pulldown543 ( pull_down543 ) ;
  TBCLL pulldown551 ( pull_down551 ) ;
  TBCLL pulldown607 ( pull_down607 ) ;
  TBCLL pulldown615 ( pull_down615 ) ;
  TBCLL pulldown623 ( pull_down623 ) ;
  TBCLL pulldown631 ( pull_down631 ) ;
  TBCLL pulldown703 ( pull_down703 ) ;
  TBCLL pulldown711 ( pull_down711 ) ;
  TBCLL pulldown288 ( pull_down288 ) ;
  TBCLL pulldown296 ( pull_down296 ) ;
  TBCLL pulldown368 ( pull_down368 ) ;
  TBCLL pulldown376 ( pull_down376 ) ;
  TBCLL pulldown384 ( pull_down384 ) ;
  TBCLL pulldown392 ( pull_down392 ) ;
  TBCLL pulldown448 ( pull_down448 ) ;
  TBCLL pulldown456 ( pull_down456 ) ;
  TBCLL pulldown464 ( pull_down464 ) ;
  TBCLL pulldown472 ( pull_down472 ) ;
  TBCLL pulldown480 ( pull_down480 ) ;
  TBCLL pulldown528 ( pull_down528 ) ;
  TBCLL pulldown536 ( pull_down536 ) ;
  TBCLL pulldown544 ( pull_down544 ) ;
  TBCLL pulldown552 ( pull_down552 ) ;
  TBCLL pulldown560 ( pull_down560 ) ;
  TBCLL pulldown608 ( pull_down608 ) ;
  TBCLL pulldown616 ( pull_down616 ) ;
  TBCLL pulldown624 ( pull_down624 ) ;
  TBCLL pulldown632 ( pull_down632 ) ;
  TBCLL pulldown640 ( pull_down640 ) ;
  TBCLL pulldown704 ( pull_down704 ) ;
  TBCLL pulldown712 ( pull_down712 ) ;
  TBCLL pulldown720 ( pull_down720 ) ;
  TBCLL pulldown289 ( pull_down289 ) ;
  TBCLL pulldown297 ( pull_down297 ) ;
  TBCLL pulldown369 ( pull_down369 ) ;
  TBCLL pulldown377 ( pull_down377 ) ;
  TBCLL pulldown385 ( pull_down385 ) ;
  TBCLL pulldown393 ( pull_down393 ) ;
  TBCLL pulldown449 ( pull_down449 ) ;
  TBCLL pulldown457 ( pull_down457 ) ;
  TBCLL pulldown465 ( pull_down465 ) ;
  TBCLL pulldown473 ( pull_down473 ) ;
  TBCLL pulldown481 ( pull_down481 ) ;
  TBCLL pulldown529 ( pull_down529 ) ;
  TBCLL pulldown537 ( pull_down537 ) ;
  TBCLL pulldown545 ( pull_down545 ) ;
  TBCLL pulldown553 ( pull_down553 ) ;
  TBCLL pulldown561 ( pull_down561 ) ;
  TBCLL pulldown609 ( pull_down609 ) ;
  TBCLL pulldown617 ( pull_down617 ) ;
  TBCLL pulldown625 ( pull_down625 ) ;
  TBCLL pulldown633 ( pull_down633 ) ;
  TBCLL pulldown641 ( pull_down641 ) ;
  TBCLL pulldown705 ( pull_down705 ) ;
  TBCLL pulldown713 ( pull_down713 ) ;
  TBCLL pulldown721 ( pull_down721 ) ;
  TBCLL pulldown298 ( pull_down298 ) ;
  TBCLL pulldown378 ( pull_down378 ) ;
  TBCLL pulldown386 ( pull_down386 ) ;
  TBCLL pulldown394 ( pull_down394 ) ;
  TBCLL pulldown458 ( pull_down458 ) ;
  TBCLL pulldown466 ( pull_down466 ) ;
  TBCLL pulldown474 ( pull_down474 ) ;
  TBCLL pulldown482 ( pull_down482 ) ;
  TBCLL pulldown490 ( pull_down490 ) ;
  TBCLL pulldown538 ( pull_down538 ) ;
  TBCLL pulldown546 ( pull_down546 ) ;
  TBCLL pulldown554 ( pull_down554 ) ;
  TBCLL pulldown562 ( pull_down562 ) ;
  TBCLL pulldown570 ( pull_down570 ) ;
  TBCLL pulldown618 ( pull_down618 ) ;
  TBCLL pulldown626 ( pull_down626 ) ;
  TBCLL pulldown634 ( pull_down634 ) ;
  TBCLL pulldown642 ( pull_down642 ) ;
  TBCLL pulldown650 ( pull_down650 ) ;
  TBCLL pulldown706 ( pull_down706 ) ;
  TBCLL pulldown714 ( pull_down714 ) ;
  TBCLL pulldown722 ( pull_down722 ) ;
  TBCLL pulldown730 ( pull_down730 ) ;
  TBCLL pulldown299 ( pull_down299 ) ;
  TBCLL pulldown379 ( pull_down379 ) ;
  TBCLL pulldown387 ( pull_down387 ) ;
  TBCLL pulldown395 ( pull_down395 ) ;
  TBCLL pulldown459 ( pull_down459 ) ;
  TBCLL pulldown467 ( pull_down467 ) ;
  TBCLL pulldown475 ( pull_down475 ) ;
  TBCLL pulldown483 ( pull_down483 ) ;
  TBCLL pulldown491 ( pull_down491 ) ;
  TBCLL pulldown539 ( pull_down539 ) ;
  TBCLL pulldown547 ( pull_down547 ) ;
  TBCLL pulldown555 ( pull_down555 ) ;
  TBCLL pulldown563 ( pull_down563 ) ;
  TBCLL pulldown571 ( pull_down571 ) ;
  TBCLL pulldown619 ( pull_down619 ) ;
  TBCLL pulldown627 ( pull_down627 ) ;
  TBCLL pulldown635 ( pull_down635 ) ;
  TBCLL pulldown643 ( pull_down643 ) ;
  TBCLL pulldown651 ( pull_down651 ) ;
  TBCLL pulldown707 ( pull_down707 ) ;
  TBCLL pulldown715 ( pull_down715 ) ;
  TBCLL pulldown723 ( pull_down723 ) ;
  TBCLL pulldown731 ( pull_down731 ) ;
  TBCLL pulldown388 ( pull_down388 ) ;
  TBCLL pulldown396 ( pull_down396 ) ;
  TBCLL pulldown468 ( pull_down468 ) ;
  TBCLL pulldown476 ( pull_down476 ) ;
  TBCLL pulldown484 ( pull_down484 ) ;
  TBCLL pulldown492 ( pull_down492 ) ;
  TBCLL pulldown548 ( pull_down548 ) ;
  TBCLL pulldown556 ( pull_down556 ) ;
  TBCLL pulldown564 ( pull_down564 ) ;
  TBCLL pulldown572 ( pull_down572 ) ;
  TBCLL pulldown580 ( pull_down580 ) ;
  TBCLL pulldown628 ( pull_down628 ) ;
  TBCLL pulldown636 ( pull_down636 ) ;
  TBCLL pulldown644 ( pull_down644 ) ;
  TBCLL pulldown652 ( pull_down652 ) ;
  TBCLL pulldown660 ( pull_down660 ) ;
  TBCLL pulldown708 ( pull_down708 ) ;
  TBCLL pulldown716 ( pull_down716 ) ;
  TBCLL pulldown724 ( pull_down724 ) ;
  TBCLL pulldown732 ( pull_down732 ) ;
  TBCLL pulldown740 ( pull_down740 ) ;
  TBCLL pulldown389 ( pull_down389 ) ;
  TBCLL pulldown397 ( pull_down397 ) ;
  TBCLL pulldown469 ( pull_down469 ) ;
  TBCLL pulldown477 ( pull_down477 ) ;
  TBCLL pulldown485 ( pull_down485 ) ;
  TBCLL pulldown493 ( pull_down493 ) ;
  TBCLL pulldown549 ( pull_down549 ) ;
  TBCLL pulldown557 ( pull_down557 ) ;
  TBCLL pulldown565 ( pull_down565 ) ;
  TBCLL pulldown573 ( pull_down573 ) ;
  TBCLL pulldown581 ( pull_down581 ) ;
  TBCLL pulldown629 ( pull_down629 ) ;
  TBCLL pulldown637 ( pull_down637 ) ;
  TBCLL pulldown645 ( pull_down645 ) ;
  TBCLL pulldown653 ( pull_down653 ) ;
  TBCLL pulldown661 ( pull_down661 ) ;
  TBCLL pulldown709 ( pull_down709 ) ;
  TBCLL pulldown717 ( pull_down717 ) ;
  TBCLL pulldown725 ( pull_down725 ) ;
  TBCLL pulldown733 ( pull_down733 ) ;
  TBCLL pulldown741 ( pull_down741 ) ;
  TBCLL pulldown398 ( pull_down398 ) ;
  TBCLL pulldown478 ( pull_down478 ) ;
  TBCLL pulldown486 ( pull_down486 ) ;
  TBCLL pulldown494 ( pull_down494 ) ;
  TBCLL pulldown558 ( pull_down558 ) ;
  TBCLL pulldown566 ( pull_down566 ) ;
  TBCLL pulldown574 ( pull_down574 ) ;
  TBCLL pulldown582 ( pull_down582 ) ;
  TBCLL pulldown590 ( pull_down590 ) ;
  TBCLL pulldown638 ( pull_down638 ) ;
  TBCLL pulldown646 ( pull_down646 ) ;
  TBCLL pulldown654 ( pull_down654 ) ;
  TBCLL pulldown662 ( pull_down662 ) ;
  TBCLL pulldown670 ( pull_down670 ) ;
  TBCLL pulldown718 ( pull_down718 ) ;
  TBCLL pulldown726 ( pull_down726 ) ;
  TBCLL pulldown734 ( pull_down734 ) ;
  TBCLL pulldown742 ( pull_down742 ) ;
  TBCLL pulldown399 ( pull_down399 ) ;
  TBCLL pulldown479 ( pull_down479 ) ;
  TBCLL pulldown487 ( pull_down487 ) ;
  TBCLL pulldown495 ( pull_down495 ) ;
  TBCLL pulldown559 ( pull_down559 ) ;
  TBCLL pulldown567 ( pull_down567 ) ;
  TBCLL pulldown575 ( pull_down575 ) ;
  TBCLL pulldown583 ( pull_down583 ) ;
  TBCLL pulldown591 ( pull_down591 ) ;
  TBCLL pulldown639 ( pull_down639 ) ;
  TBCLL pulldown647 ( pull_down647 ) ;
  TBCLL pulldown655 ( pull_down655 ) ;
  TBCLL pulldown663 ( pull_down663 ) ;
  TBCLL pulldown671 ( pull_down671 ) ;
  TBCLL pulldown719 ( pull_down719 ) ;
  TBCLL pulldown727 ( pull_down727 ) ;
  TBCLL pulldown735 ( pull_down735 ) ;
  TBCLL pulldown743 ( pull_down743 ) ;
  TBCLL pulldown488 ( pull_down488 ) ;
  TBCLL pulldown496 ( pull_down496 ) ;
  TBCLL pulldown568 ( pull_down568 ) ;
  TBCLL pulldown576 ( pull_down576 ) ;
  TBCLL pulldown584 ( pull_down584 ) ;
  TBCLL pulldown592 ( pull_down592 ) ;
  TBCLL pulldown648 ( pull_down648 ) ;
  TBCLL pulldown656 ( pull_down656 ) ;
  TBCLL pulldown664 ( pull_down664 ) ;
  TBCLL pulldown672 ( pull_down672 ) ;
  TBCLL pulldown680 ( pull_down680 ) ;
  TBCLL pulldown728 ( pull_down728 ) ;
  TBCLL pulldown736 ( pull_down736 ) ;
  TBCLL pulldown744 ( pull_down744 ) ;
  TBCLL pulldown489 ( pull_down489 ) ;
  TBCLL pulldown497 ( pull_down497 ) ;
  TBCLL pulldown569 ( pull_down569 ) ;
  TBCLL pulldown577 ( pull_down577 ) ;
  TBCLL pulldown585 ( pull_down585 ) ;
  TBCLL pulldown593 ( pull_down593 ) ;
  TBCLL pulldown649 ( pull_down649 ) ;
  TBCLL pulldown657 ( pull_down657 ) ;
  TBCLL pulldown665 ( pull_down665 ) ;
  TBCLL pulldown673 ( pull_down673 ) ;
  TBCLL pulldown681 ( pull_down681 ) ;
  TBCLL pulldown729 ( pull_down729 ) ;
  TBCLL pulldown737 ( pull_down737 ) ;
  TBCLL pulldown745 ( pull_down745 ) ;
  TBCLL pulldown498 ( pull_down498 ) ;
  TBCLL pulldown578 ( pull_down578 ) ;
  TBCLL pulldown586 ( pull_down586 ) ;
  TBCLL pulldown594 ( pull_down594 ) ;
  TBCLL pulldown658 ( pull_down658 ) ;
  TBCLL pulldown666 ( pull_down666 ) ;
  TBCLL pulldown674 ( pull_down674 ) ;
  TBCLL pulldown682 ( pull_down682 ) ;
  TBCLL pulldown690 ( pull_down690 ) ;
  TBCLL pulldown738 ( pull_down738 ) ;
  TBCLL pulldown746 ( pull_down746 ) ;
  TBCLL pulldown499 ( pull_down499 ) ;
  TBCLL pulldown579 ( pull_down579 ) ;
  TBCLL pulldown587 ( pull_down587 ) ;
  TBCLL pulldown595 ( pull_down595 ) ;
  TBCLL pulldown659 ( pull_down659 ) ;
  TBCLL pulldown667 ( pull_down667 ) ;
  TBCLL pulldown675 ( pull_down675 ) ;
  TBCLL pulldown683 ( pull_down683 ) ;
  TBCLL pulldown691 ( pull_down691 ) ;
  TBCLL pulldown739 ( pull_down739 ) ;
  TBCLL pulldown747 ( pull_down747 ) ;
  TBCLL pulldown588 ( pull_down588 ) ;
  TBCLL pulldown596 ( pull_down596 ) ;
  TBCLL pulldown668 ( pull_down668 ) ;
  TBCLL pulldown676 ( pull_down676 ) ;
  TBCLL pulldown684 ( pull_down684 ) ;
  TBCLL pulldown692 ( pull_down692 ) ;
  TBCLL pulldown589 ( pull_down589 ) ;
  TBCLL pulldown597 ( pull_down597 ) ;
  TBCLL pulldown669 ( pull_down669 ) ;
  TBCLL pulldown677 ( pull_down677 ) ;
  TBCLL pulldown685 ( pull_down685 ) ;
  TBCLL pulldown693 ( pull_down693 ) ;
  TBCLL pulldown598 ( pull_down598 ) ;
  TBCLL pulldown678 ( pull_down678 ) ;
  TBCLL pulldown686 ( pull_down686 ) ;
  TBCLL pulldown694 ( pull_down694 ) ;
  TBCLL pulldown599 ( pull_down599 ) ;
  TBCLL pulldown679 ( pull_down679 ) ;
  TBCLL pulldown687 ( pull_down687 ) ;
  TBCLL pulldown695 ( pull_down695 ) ;
  TBCLL pulldown688 ( pull_down688 ) ;
  TBCLL pulldown696 ( pull_down696 ) ;
  TBCLL pulldown689 ( pull_down689 ) ;
  TBCLL pulldown697 ( pull_down697 ) ;
  TBCLL pulldown698 ( pull_down698 ) ;
  TBCLL pulldown699 ( pull_down699 ) ;
  TBCLH pullup0 ( pull_up0 ) ;
  TBCLH pullup1 ( pull_up1 ) ;
  TBCLH pullup2 ( pull_up2 ) ;
  TBCLH pullup3 ( pull_up3 ) ;
  TBCLH pullup4 ( pull_up4 ) ;

  // Refer to /proj/78k0r_11/78k0r_kx4/_ice/_make_chip/_chiptop/_library/chiptop_045.v
  chiptop chiptop (
    .MDRRAM15 ( MDRRAM15 ) ,.MDRRAM14 ( MDRRAM14 ) ,.MDRRAM13 ( MDRRAM13 )
     ,.MDRRAM12 ( MDRRAM12 ) ,.MDRRAM11 ( MDRRAM11 ) ,.MDRRAM10 ( MDRRAM10 )
     ,.MDRRAM9 ( MDRRAM9 ) ,.MDRRAM8 ( MDRRAM8 ) ,.MDRRAM7 ( MDRRAM7 )
     ,.MDRRAM6 ( MDRRAM6 ) ,.MDRRAM5 ( MDRRAM5 ) ,.MDRRAM4 ( MDRRAM4 )
     ,.MDRRAM3 ( MDRRAM3 ) ,.MDRRAM2 ( MDRRAM2 ) ,.MDRRAM1 ( MDRRAM1 )
     ,.MDRRAM0 ( MDRRAM0 ) ,.A19 ( A19 ) ,.A18 ( A18 ) ,.A17 ( A17 ) ,.A16 ( A16 )
     ,.A15 ( A15 ) ,.A14 ( A14 ) ,.A13 ( A13 ) ,.A12 ( A12 ) ,.A11 ( A11 )
     ,.A10 ( A10 ) ,.A9 ( A9 ) ,.A8 ( A8 ) ,.A7 ( A7 ) ,.A6 ( A6 ) ,.A5 ( A5 )
     ,.A4 ( A4 ) ,.A3 ( A3 ) ,.A2 ( A2 ) ,.CE0 ( CE0 ) ,.DA4 ( DA4 ) ,.AF6 ( AF6 )
     ,.CE1 ( CE1 ) ,.DA5 ( DA5 ) ,.AF7 ( AF7 ) ,.SELRO1 ( SELRO1 ) ,.CLKSEL1 ( CLKSEL1 )
     ,.EXA ( EXA ) ,.BFA ( BFA ) ,.ICETMSPMD ( ICETMSPMD ) ,.ICETMBTSEL ( ICETMBTSEL )
     ,.BRSAM ( BRSAM ) ,.PID31 ( CIBPID31 ) ,.PID23 ( CIBPID23 ) ,.PID15 ( CIBPID15 )
     ,.RO111 ( RO111 ) ,.RO031 ( RO031 ) ,.RO023 ( RO023 ) ,.RO015 ( RO015 )
     ,.PID30 ( CIBPID30 ) ,.PID22 ( CIBPID22 ) ,.PID14 ( CIBPID14 ) ,.RO110 ( RO110 )
     ,.RO030 ( RO030 ) ,.RO022 ( RO022 ) ,.RO014 ( RO014 ) ,.PID29 ( CIBPID29 )
     ,.RO133 ( RO133 ) ,.RO125 ( RO125 ) ,.RO117 ( RO117 ) ,.RO037 ( RO037 )
     ,.RO029 ( RO029 ) ,.PID28 ( CIBPID28 ) ,.RO132 ( RO132 ) ,.RO124 ( RO124 )
     ,.RO116 ( RO116 ) ,.RO036 ( RO036 ) ,.RO028 ( RO028 ) ,.PID27 ( CIBPID27 )
     ,.PID19 ( CIBPID19 ) ,.RO131 ( RO131 ) ,.RO123 ( RO123 ) ,.RO115 ( RO115 )
     ,.RO035 ( RO035 ) ,.RO027 ( RO027 ) ,.RO019 ( RO019 ) ,.PID26 ( CIBPID26 )
     ,.PID18 ( CIBPID18 ) ,.RO130 ( RO130 ) ,.RO122 ( RO122 ) ,.RO114 ( RO114 )
     ,.RO034 ( RO034 ) ,.RO026 ( RO026 ) ,.RO018 ( RO018 ) ,.PID25 ( CIBPID25 )
     ,.PID17 ( CIBPID17 ) ,.RO121 ( RO121 ) ,.RO113 ( RO113 ) ,.RO033 ( RO033 )
     ,.RO025 ( RO025 ) ,.RO017 ( RO017 ) ,.PID24 ( CIBPID24 ) ,.PID16 ( CIBPID16 )
     ,.RO120 ( RO120 ) ,.RO112 ( RO112 ) ,.RO032 ( RO032 ) ,.RO024 ( RO024 )
     ,.RO016 ( RO016 ) ,.PID21 ( CIBPID21 ) ,.PID13 ( CIBPID13 ) ,.RO021 ( RO021 )
     ,.RO013 ( RO013 ) ,.PID20 ( CIBPID20 ) ,.PID12 ( CIBPID12 ) ,.RO020 ( RO020 )
     ,.RO012 ( RO012 ) ,.CPURD ( CPURD ) ,.PID11 ( CIBPID11 ) ,.RO011 ( RO011 )
     ,.PID10 ( CIBPID10 ) ,.RO010 ( RO010 ) ,.PID9 ( CIBPID9 ) ,.RO17 ( RO17 )
     ,.RO09 ( RO09 ) ,.PID8 ( CIBPID8 ) ,.RO16 ( RO16 ) ,.RO08 ( RO08 )
     ,.PID7 ( CIBPID7 ) ,.RO15 ( RO15 ) ,.RO07 ( RO07 ) ,.PID6 ( CIBPID6 )
     ,.RO14 ( RO14 ) ,.RO06 ( RO06 ) ,.PID5 ( CIBPID5 ) ,.RO13 ( RO13 )
     ,.RO05 ( RO05 ) ,.PID4 ( CIBPID4 ) ,.RO12 ( RO12 ) ,.RO04 ( RO04 )
     ,.PID3 ( CIBPID3 ) ,.RO11 ( RO11 ) ,.RO03 ( RO03 ) ,.MDW9 ( MDW9 )
     ,.PID2 ( CIBPID2 ) ,.RO10 ( RO10 ) ,.RO02 ( RO02 ) ,.MDW8 ( MDW8 )
     ,.PID1 ( CIBPID1 ) ,.RO01 ( RO01 ) ,.MDW7 ( MDW7 ) ,.PID0 ( CIBPID0 )
     ,.RO00 ( RO00 ) ,.MDW6 ( MDW6 ) ,.RO137 ( RO137 ) ,.RO129 ( RO129 )
     ,.EXMA3 ( EXMA3 ) ,.FLSPM ( FLSPM ) ,.RO136 ( RO136 ) ,.RO128 ( RO128 )
     ,.EXMA2 ( EXMA2 ) ,.RO135 ( RO135 ) ,.RO127 ( RO127 ) ,.RO119 ( RO119 )
     ,.EXMA1 ( EXMA1 ) ,.RO134 ( RO134 ) ,.RO126 ( RO126 ) ,.RO118 ( RO118 )
     ,.EXMA0 ( EXMA0 ) ,.RO19 ( RO19 ) ,.RO18 ( RO18 ) ,.DCE0 ( DCE0 )
     ,.DCLKSEL1 ( DCLKSEL1 ) ,.DRDCLKC1 ( DRDCLKC1 ) ,.DA13 ( DA13 ) ,.AF17 ( AF17 )
     ,.DA12 ( DA12 ) ,.AF16 ( AF16 ) ,.DA11 ( DA11 ) ,.AF15 ( AF15 ) ,.DA10 ( DA10 )
     ,.AF14 ( AF14 ) ,.DA9 ( DA9 ) ,.DA8 ( DA8 ) ,.DA7 ( DA7 ) ,.AF9 ( AF9 )
     ,.DA6 ( DA6 ) ,.AF8 ( AF8 ) ,.DA3 ( DA3 ) ,.AF5 ( AF5 ) ,.DA2 ( DA2 )
     ,.AF4 ( AF4 ) ,.DA1 ( DA1 ) ,.AF3 ( AF3 ) ,.DA0 ( DA0 ) ,.AF2 ( AF2 )
     ,.DRO00 ( DRO00 ) ,.DRO01 ( DRO01 ) ,.DRO02 ( DRO02 ) ,.DRO03 ( DRO03 )
     ,.DRO04 ( DRO04 ) ,.DRO05 ( DRO05 ) ,.DRO06 ( DRO06 ) ,.DRO07 ( DRO07 )
     ,.DRO08 ( DRO08 ) ,.DRO09 ( DRO09 ) ,.DRO010 ( DRO010 ) ,.DRO011 ( DRO011 )
     ,.SLFLASH ( SLFLASH ) ,.WAITFL2 ( WAITFL2 ) ,.SVI ( SVI ) ,.SVVCOUT7 ( SVVCOUT7 )
     ,.SVVCOUT6 ( SVVCOUT6 ) ,.SVVCOUT5 ( SVVCOUT5 ) ,.SVVCOUT4 ( SVVCOUT4 )
     ,.SVVCOUT3 ( SVVCOUT3 ) ,.SVVCOUT2 ( SVVCOUT2 ) ,.SVVCOUT1 ( SVVCOUT1 )
     ,.SVVCOUT0 ( SVVCOUT0 ) ,.SVINTACK ( SVINTACK ) ,.SOFTBRK ( SOFTBRK )
     ,.ICEMSKNMI ( ICEMSKNMI ) ,.ICEMSKDBG ( ICEMSKDBG ) ,.STAGEADR1 ( STAGEADR1 )
     ,.STAGEADR0 ( STAGEADR0 ) ,.PREFIX ( PREFIX ) ,.SKIPEXE ( SKIPEXE )
     ,.PCWAITF ( PCWAITF ) ,.CPUMASK ( CPUMASK ) ,.CPUPID1 ( CPUPID1 )
     ,.CPUMISAL ( CPUMISAL ) ,.FLREAD ( FLREAD ) ,.IMDR10 ( IMDR10 ) ,.FLREADB3 ( FLREADB3 )
     ,.FLREADB2 ( FLREADB2 ) ,.FLREADB1 ( FLREADB1 ) ,.FLREADB0 ( FLREADB0 )
     ,.FCHRAM ( FCHRAM ) ,.SLMEM ( SLMEM ) ,.SLEXM ( SLEXM ) ,.SLBMEM ( SLBMEM )
     ,.SPDEC ( SPDEC ) ,.SPINC ( SPINC ) ,.SPREL ( SPREL ) ,.IDPOP ( IDPOP )
     ,.MDW10 ( MDW10 ) ,.IMDR2 ( IMDR2 ) ,.CPUWR ( CPUWR ) ,.WDOP ( WDOP )
     ,.ICEWAITMEM ( ICEWAITMEM ) ,.DMAACK ( DMAACK ) ,.HLTST ( HLTST )
     ,.STPST ( STPST ) ,.INTACK ( INTACK ) ,.OCDWAIT ( OCDWAIT ) ,.SVMOD ( SVMOD )
     ,.SVMODF ( SVMODF ) ,.ALT1 ( ALT1 ) ,.DW21 ( DW21 ) ,.DW13 ( DW13 )
     ,.DRDCLK ( DRDCLK ) ,.SLDFLASH ( SLDFLASH ) ,.ICECSGREGU ( ICECSGREGU )
     ,.ICEIFA4 ( ICEIFA4 ) ,.ICEIFA3 ( ICEIFA3 ) ,.ICEIFA2 ( ICEIFA2 )
     ,.ICEDO31 ( ICEDO31 ) ,.ICEDO23 ( ICEDO23 ) ,.ICEDO15 ( ICEDO15 )
     ,.ICEDO30 ( ICEDO30 ) ,.ICEDO22 ( ICEDO22 ) ,.ICEDO14 ( ICEDO14 )
     ,.ICEDO29 ( ICEDO29 ) ,.ICEDO28 ( ICEDO28 ) ,.ICEDO27 ( ICEDO27 )
     ,.ICEDO19 ( ICEDO19 ) ,.ICEDO26 ( ICEDO26 ) ,.ICEDO18 ( ICEDO18 )
     ,.ICEDO25 ( ICEDO25 ) ,.ICEDO17 ( ICEDO17 ) ,.ICEDO24 ( ICEDO24 )
     ,.ICEDO16 ( ICEDO16 ) ,.ICEDO21 ( ICEDO21 ) ,.ICEDO13 ( ICEDO13 )
     ,.ICEDO20 ( ICEDO20 ) ,.ICEDO12 ( ICEDO12 ) ,.P74PUON ( P74PUON )
     ,.ICEDO11 ( ICEDO11 ) ,.ICEDO10 ( ICEDO10 ) ,.ICEDO9 ( ICEDO9 ) ,.ICEDO8 ( ICEDO8 )
     ,.ICEDO7 ( ICEDO7 ) ,.ICEDO6 ( ICEDO6 ) ,.ICEDO5 ( ICEDO5 ) ,.ICEDO4 ( ICEDO4 )
     ,.ICEDO3 ( ICEDO3 ) ,.ICEDO2 ( ICEDO2 ) ,.ICEDO1 ( ICEDO1 ) ,.ICEDO0 ( ICEDO0 )
     ,.PA19 ( PA19 ) ,.PC11 ( PC11 ) ,.PA18 ( PA18 ) ,.PC10 ( PC10 ) ,.PA17 ( PA17 )
     ,.PA16 ( PA16 ) ,.PA15 ( PA15 ) ,.PA14 ( PA14 ) ,.PA13 ( PA13 ) ,.DW37 ( DW37 )
     ,.DW29 ( DW29 ) ,.PA12 ( PA12 ) ,.DW36 ( DW36 ) ,.DW28 ( DW28 ) ,.PA11 ( PA11 )
     ,.DW35 ( DW35 ) ,.DW27 ( DW27 ) ,.DW19 ( DW19 ) ,.PA10 ( PA10 ) ,.DW34 ( DW34 )
     ,.DW26 ( DW26 ) ,.DW18 ( DW18 ) ,.PA9 ( PA9 ) ,.PC5 ( PC5 ) ,.PA8 ( PA8 )
     ,.PC4 ( PC4 ) ,.PA7 ( PA7 ) ,.PC3 ( PC3 ) ,.PA6 ( PA6 ) ,.PC2 ( PC2 )
     ,.PA5 ( PA5 ) ,.PC1 ( PC1 ) ,.DW9 ( DW9 ) ,.PA4 ( PA4 ) ,.PC0 ( PC0 )
     ,.DW8 ( DW8 ) ,.PA3 ( PA3 ) ,.DW7 ( DW7 ) ,.DIS ( DIS ) ,.PA2 ( PA2 )
     ,.DW6 ( DW6 ) ,.PC19 ( PC19 ) ,.PC18 ( PC18 ) ,.PC17 ( PC17 ) ,.PC16 ( PC16 )
     ,.PC15 ( PC15 ) ,.PC14 ( PC14 ) ,.PC13 ( PC13 ) ,.PC12 ( PC12 ) ,.PC9 ( PC9 )
     ,.PC8 ( PC8 ) ,.PC7 ( PC7 ) ,.PC6 ( PC6 ) ,.IDADR31 ( IDADR31 ) ,.IDADR23 ( IDADR23 )
     ,.IDADR15 ( IDADR15 ) ,.ICEDI19 ( ICEDI19 ) ,.ICEDI27 ( ICEDI27 )
     ,.IDADR30 ( IDADR30 ) ,.IDADR22 ( IDADR22 ) ,.IDADR14 ( IDADR14 )
     ,.ICEDI18 ( ICEDI18 ) ,.ICEDI26 ( ICEDI26 ) ,.IDADR29 ( IDADR29 )
     ,.IDADR28 ( IDADR28 ) ,.IDADR27 ( IDADR27 ) ,.IDADR19 ( IDADR19 )
     ,.IDADR26 ( IDADR26 ) ,.IDADR18 ( IDADR18 ) ,.IDADR25 ( IDADR25 )
     ,.IDADR17 ( IDADR17 ) ,.ICEDI29 ( ICEDI29 ) ,.IDADR24 ( IDADR24 )
     ,.IDADR16 ( IDADR16 ) ,.ICEDI28 ( ICEDI28 ) ,.P73PUON ( P73PUON )
     ,.IDADR21 ( IDADR21 ) ,.IDADR13 ( IDADR13 ) ,.ICEDI17 ( ICEDI17 )
     ,.ICEDI25 ( ICEDI25 ) ,.IDADR20 ( IDADR20 ) ,.IDADR12 ( IDADR12 )
     ,.ICEDI16 ( ICEDI16 ) ,.ICEDI24 ( ICEDI24 ) ,.IDADR11 ( IDADR11 )
     ,.ICEDI15 ( ICEDI15 ) ,.ICEDI23 ( ICEDI23 ) ,.ICEDI31 ( ICEDI31 )
     ,.IDADR10 ( IDADR10 ) ,.ICEDI14 ( ICEDI14 ) ,.ICEDI22 ( ICEDI22 )
     ,.ICEDI30 ( ICEDI30 ) ,.IDADR9 ( IDADR9 ) ,.IDADR8 ( IDADR8 ) ,.IDADR7 ( IDADR7 )
     ,.ICEDI9 ( ICEDI9 ) ,.IDADR6 ( IDADR6 ) ,.ICEDI8 ( ICEDI8 ) ,.IDADR5 ( IDADR5 )
     ,.ICEDI7 ( ICEDI7 ) ,.IDADR4 ( IDADR4 ) ,.ICEDI6 ( ICEDI6 ) ,.IDADR3 ( IDADR3 )
     ,.ICEDI5 ( ICEDI5 ) ,.IDADR2 ( IDADR2 ) ,.ICEDI4 ( ICEDI4 ) ,.IDADR1 ( IDADR1 )
     ,.ICEDI3 ( ICEDI3 ) ,.IDADR0 ( IDADR0 ) ,.ICEDI2 ( ICEDI2 ) ,.MA15 ( MA15 )
     ,.MA14 ( MA14 ) ,.MA13 ( MA13 ) ,.MA12 ( MA12 ) ,.BEU2 ( BEU2 ) ,.MA11 ( MA11 )
     ,.BEU1 ( BEU1 ) ,.MA10 ( MA10 ) ,.BEU0 ( BEU0 ) ,.MA9 ( MA9 ) ,.DW1 ( DW1 )
     ,.MA8 ( MA8 ) ,.DW0 ( DW0 ) ,.MA7 ( MA7 ) ,.MA6 ( MA6 ) ,.MA5 ( MA5 )
     ,.MA4 ( MA4 ) ,.MA3 ( MA3 ) ,.MA2 ( MA2 ) ,.CER ( CER ) ,.MA1 ( MA1 )
     ,.MA0 ( MA0 ) ,.MDW15 ( MDW15 ) ,.IMDR7 ( IMDR7 ) ,.MDW14 ( MDW14 )
     ,.IMDR6 ( IMDR6 ) ,.MDW13 ( MDW13 ) ,.IMDR5 ( IMDR5 ) ,.MDW12 ( MDW12 )
     ,.IMDR4 ( IMDR4 ) ,.MDW11 ( MDW11 ) ,.IMDR3 ( IMDR3 ) ,.MDW5 ( MDW5 )
     ,.MDW4 ( MDW4 ) ,.MDW3 ( MDW3 ) ,.MDW2 ( MDW2 ) ,.MDW1 ( MDW1 ) ,.MDW0 ( MDW0 )
     ,.EXCH ( EXCH ) ,.IMDR15 ( IMDR15 ) ,.IMDR14 ( IMDR14 ) ,.IMDR13 ( IMDR13 )
     ,.IMDR12 ( IMDR12 ) ,.IMDR11 ( IMDR11 ) ,.IMDR9 ( IMDR9 ) ,.IMDR8 ( IMDR8 )
     ,.IMDR1 ( IMDR1 ) ,.IMDR0 ( IMDR0 ) ,.CPUPID31 ( CPUPID31 ) ,.CPUPID23 ( CPUPID23 )
     ,.CPUPID15 ( CPUPID15 ) ,.CPUPID30 ( CPUPID30 ) ,.CPUPID22 ( CPUPID22 )
     ,.CPUPID14 ( CPUPID14 ) ,.CPUPID29 ( CPUPID29 ) ,.CPUPID28 ( CPUPID28 )
     ,.CPUPID27 ( CPUPID27 ) ,.CPUPID19 ( CPUPID19 ) ,.CPUPID26 ( CPUPID26 )
     ,.CPUPID18 ( CPUPID18 ) ,.CPUPID25 ( CPUPID25 ) ,.CPUPID17 ( CPUPID17 )
     ,.CPUPID24 ( CPUPID24 ) ,.CPUPID16 ( CPUPID16 ) ,.CPUPID21 ( CPUPID21 )
     ,.CPUPID13 ( CPUPID13 ) ,.CPUPID20 ( CPUPID20 ) ,.CPUPID12 ( CPUPID12 )
     ,.CPUPID11 ( CPUPID11 ) ,.CPUPID10 ( CPUPID10 ) ,.CPUPID9 ( CPUPID9 )
     ,.CPUPID8 ( CPUPID8 ) ,.CPUPID7 ( CPUPID7 ) ,.CPUPID6 ( CPUPID6 )
     ,.CPUPID5 ( CPUPID5 ) ,.CPUPID4 ( CPUPID4 ) ,.CPUPID3 ( CPUPID3 )
     ,.CPUPID2 ( CPUPID2 ) ,.CPUPID0 ( CPUPID0 ) ,.FLSIZE3 ( FLSIZE3 )
     ,.FLSIZE2 ( FLSIZE2 ) ,.FLSIZE1 ( FLSIZE1 ) ,.FLSIZE0 ( FLSIZE0 )
     ,.RAMSIZE7 ( RAMSIZE7 ) ,.RAMSIZE6 ( RAMSIZE6 ) ,.RAMSIZE5 ( RAMSIZE5 )
     ,.RAMSIZE4 ( RAMSIZE4 ) ,.RAMSIZE3 ( RAMSIZE3 ) ,.RAMSIZE2 ( RAMSIZE2 )
     ,.RAMSIZE1 ( RAMSIZE1 ) ,.RAMSIZE0 ( RAMSIZE0 ) ,.BFSIZE3 ( BFSIZE3 )
     ,.BFSIZE2 ( BFSIZE2 ) ,.BFSIZE1 ( BFSIZE1 ) ,.BFSIZE0 ( BFSIZE0 )
     ,.BMSIZE3 ( BMSIZE3 ) ,.BMSIZE2 ( BMSIZE2 ) ,.BMSIZE1 ( BMSIZE1 )
     ,.BMSIZE0 ( BMSIZE0 ) ,.DFSIZE1 ( DFSIZE1 ) ,.DFSIZE0 ( DFSIZE0 )
     ,.ICEMKLVI ( ICEMKLVI ) ,.ICEMKWDT ( ICEMKWDT ) ,.RESETB ( RESETB )
     ,.RESB ( RESB ) ,.FCLKRT ( FCLK_ICE ) ,.FCLK1 ( FCLK1 ) ,.FCLK2 ( FCLK2 )
     ,.DW33 ( DW33 ) ,.DW25 ( DW25 ) ,.DW17 ( DW17 ) ,.DDIS ( DDIS ) ,.DW32 ( DW32 )
     ,.DW24 ( DW24 ) ,.DW16 ( DW16 ) ,.DW31 ( DW31 ) ,.DW23 ( DW23 ) ,.DW15 ( DW15 )
     ,.DW30 ( DW30 ) ,.DW22 ( DW22 ) ,.DW14 ( DW14 ) ,.DW20 ( DW20 ) ,.DW12 ( DW12 )
     ,.DW11 ( DW11 ) ,.DW10 ( DW10 ) ,.DW5 ( DW5 ) ,.DW4 ( DW4 ) ,.DW3 ( DW3 )
     ,.DW2 ( DW2 ) ,.TMSPMD ( TMSPMD ) ,.TMBTSEL ( TMBTSEL ) ,.BTFLG ( BTFLG )
     ,.READ ( READ ) ,.RDCLKP1 ( RDCLKP1 ) ,.SER ( SER ) ,.WED ( WED )
     ,.WWR ( WWR ) ,.MRG00 ( MRG00 ) ,.MRG01 ( MRG01 ) ,.MRG10 ( MRG10 )
     ,.MRG11 ( MRG11 ) ,.MRG12 ( MRG12 ) ,.PROGI ( PROGI ) ,.ICEFLERR ( ICEFLERR )
     ,.ICENOECC ( ICENOECC ) ,.DCER ( DCER ) ,.DSER ( DSER ) ,.DWWR ( DWWR )
     ,.DWED ( DWED ) ,.DMRG00 ( DMRG00 ) ,.DMRG01 ( DMRG01 ) ,.DMRG10 ( DMRG10 )
     ,.DMRG11 ( DMRG11 ) ,.DMRG12 ( DMRG12 ) ,.DREAD ( DREAD ) ,.AF19 ( AF19 )
     ,.AF18 ( AF18 ) ,.AF13 ( AF13 ) ,.AF12 ( AF12 ) ,.AF11 ( AF11 ) ,.AF10 ( AF10 )
     ,.AF1 ( AF1 ) ,.AF0 ( AF0 ) ,.OCDMOD ( OCDMOD ) ,.CLK60MHZ ( CLK60MHZ )
     ,.CLK30MHZ_GB ( CLK30MHZ_GB ) ,.GDRAMWR ( GDRAMWR ) ,.PSEUDOON10 ( PSEUDOON10 )
     ,.PERISVIB ( PERISVIB ) ,.PSEUDOON1 ( PSEUDOON1 ) ,.SVMODI ( SVMODI )
     ,.SVMODIPERI1 ( SVMODIPERI1 ) ,.SVMODIPERI2 ( SVMODIPERI2 ) ,.STBRELESV ( STBRELESV )
     ,.CLK30MHZ ( CLK30MHZ ) ,.LOCK48FAIL ( LOCK48FAIL ) ,.LOCK64FAIL ( LOCK64FAIL )
     ,.LOCKHROSCFAIL ( LOCKHROSCFAIL ) ,.PONRESB ( PONRESB ) ,.CPUPRCLK3 ( CPUPRCLK3 )
     ,.CPURCLK3 ( CPURCLK3 ) ,.P121 ( P121 ) ,.P122 ( P122 ) ,.CPUTMCLK ( CPUTMCLK )
     ,.CPUMCLK ( CPUMCLK ) ,.CPUTSCLK ( CPUTSCLK ) ,.CPUSCLK ( CPUSCLK )
     ,.P123 ( P123 ) ,.P124 ( P124 ) ,.POCRESB ( POCRESB ) ,.VDDLEV0 ( VDDLEV0 )
     ,.VDDLEV1 ( VDDLEV1 ) ,.VDDLEV2 ( VDDLEV2 ) ,.VDDLEV3 ( VDDLEV3 )
     ,.VDDLEV4 ( VDDLEV4 ) ,.VDDLEV5 ( VDDLEV5 ) ,.VDDLEV6 ( VDDLEV6 )
     ,.VDDLEV7 ( VDDLEV7 ) ,.USBIFWR ( USBIFWR ) ,.PSEUDOON0 ( PSEUDOON0 )
     ,.PSEUDOON8 ( PSEUDOON8 ) ,.RESINB ( RESINB ) ,.RESFB5V ( RESFB5V )
     ,.ICEDATAFLT ( PSEUDOON5 ) ,.ICEDMAFLT ( PSEUDOON6 ) ,.ICEFETCHFLT ( PSEUDOON4 )
     ,.PSEUDOTIIDER ( PSEUDOON7 ) ,.ICEMSKCKSMER ( PSEUDOON2 ) ,.PSEUDOCKSMER ( PSEUDOON3 )
     ,.SYSRSOUTB ( SYSRSOUTB ) ,.ICEWR ( ICEWR ) ,.ICEIFA0 ( ICEIFA0 )
     ,.ICEIFA1 ( ICEIFA1 ) ,.ICEIFA5 ( ICEIFA5 ) ,.ICEIFA6 ( ICEIFA6 )
     ,.ICEIFA7 ( ICEIFA7 ) ,.ICEIFA8 ( ICEIFA8 ) ,.ICEIFA9 ( ICEIFA9 )
     ,.ICEIFA10 ( ICEIFA10 ) ,.ICEIFA11 ( ICEIFA11 ) ,.ICEIFA12 ( ICEIFA12 )
     ,.ICEIFA20 ( ICEIFA20 ) ,.ICEIFA13 ( ICEIFA13 ) ,.ICEIFA21 ( ICEIFA21 )
     ,.ICEIFA14 ( ICEIFA14 ) ,.ICEIFA22 ( ICEIFA22 ) ,.ICEIFA30 ( ICEIFA30 )
     ,.ICEIFA15 ( ICEIFA15 ) ,.ICEIFA23 ( ICEIFA23 ) ,.ICEIFA31 ( ICEIFA31 )
     ,.ICEIFA16 ( ICEIFA16 ) ,.ICEIFA24 ( ICEIFA24 ) ,.ICEIFA17 ( ICEIFA17 )
     ,.ICEIFA25 ( ICEIFA25 ) ,.ICEIFA18 ( ICEIFA18 ) ,.ICEIFA26 ( ICEIFA26 )
     ,.ICEIFA19 ( ICEIFA19 ) ,.ICEIFA27 ( ICEIFA27 ) ,.ICEIFA28 ( ICEIFA28 )
     ,.ICEIFA29 ( ICEIFA29 ) ,.ICEDI0 ( ICEDI0 ) ,.ICEDI1 ( ICEDI1 ) ,.ICEDI10 ( ICEDI10 )
     ,.ICEDI11 ( ICEDI11 ) ,.ICEDI12 ( ICEDI12 ) ,.ICEDI20 ( ICEDI20 )
     ,.ICEDI13 ( ICEDI13 ) ,.ICEDI21 ( ICEDI21 ) ,.ICEDOP0 ( ICEDOP0 )
     ,.ICEDOP1 ( ICEDOP1 ) ,.ICEDOP2 ( ICEDOP2 ) ,.ICEDOP3 ( ICEDOP3 )
     ,.ICEDOP4 ( ICEDOP4 ) ,.ICEDOP5 ( ICEDOP5 ) ,.ICEDOP6 ( ICEDOP6 )
     ,.ICEDOP7 ( ICEDOP7 ) ,.ICEDOP8 ( ICEDOP8 ) ,.ICEDOP9 ( ICEDOP9 )
     ,.ICEDOP10 ( ICEDOP10 ) ,.ICEDOP11 ( ICEDOP11 ) ,.ICEDOP12 ( ICEDOP12 )
     ,.ICEDOP20 ( ICEDOP20 ) ,.ICEDOP13 ( ICEDOP13 ) ,.ICEDOP21 ( ICEDOP21 )
     ,.ICEDOP14 ( ICEDOP14 ) ,.ICEDOP22 ( ICEDOP22 ) ,.ICEDOP30 ( ICEDOP30 )
     ,.ICEDOP15 ( ICEDOP15 ) ,.ICEDOP23 ( ICEDOP23 ) ,.ICEDOP31 ( ICEDOP31 )
     ,.ICEDOP16 ( ICEDOP16 ) ,.ICEDOP24 ( ICEDOP24 ) ,.ICEDOP17 ( ICEDOP17 )
     ,.ICEDOP25 ( ICEDOP25 ) ,.ICEDOP18 ( ICEDOP18 ) ,.ICEDOP26 ( ICEDOP26 )
     ,.ICEDOP19 ( ICEDOP19 ) ,.ICEDOP27 ( ICEDOP27 ) ,.ICEDOP28 ( ICEDOP28 )
     ,.ICEDOP29 ( ICEDOP29 ) ,.STOPZ ( STOPZ ) ,.P00ENO ( P00ENO ) ,.P01ENO ( P01ENO )
     ,.P02ENO ( P02ENO ) ,.P10ENO ( P10ENO ) ,.P03ENO ( P03ENO ) ,.P11ENO ( P11ENO )
     ,.P04ENO ( P04ENO ) ,.P12ENO ( P12ENO ) ,.P20ENO ( P20ENO ) ,.P05ENO ( P05ENO )
     ,.P13ENO ( P13ENO ) ,.P21ENO ( P21ENO ) ,.P06ENO ( P06ENO ) ,.P14ENO ( P14ENO )
     ,.P22ENO ( P22ENO ) ,.P30ENO ( P30ENO ) ,.P00DOUT ( P00DOUT ) ,.P01DOUT ( P01DOUT )
     ,.P02DOUT ( P02DOUT ) ,.P10DOUT ( P10DOUT ) ,.P03DOUT ( P03DOUT )
     ,.P11DOUT ( P11DOUT ) ,.P04DOUT ( P04DOUT ) ,.P12DOUT ( P12DOUT )
     ,.P20DOUT ( P20DOUT ) ,.P05DOUT ( P05DOUT ) ,.P13DOUT ( P13DOUT )
     ,.P21DOUT ( P21DOUT ) ,.P06DOUT ( P06DOUT ) ,.P14DOUT ( P14DOUT )
     ,.P22DOUT ( P22DOUT ) ,.P30DOUT ( P30DOUT ) ,.P00ENI ( P00ENI ) ,.P01ENI ( P01ENI )
     ,.P02ENI ( P02ENI ) ,.P10ENI ( P10ENI ) ,.P03ENI ( P03ENI ) ,.P11ENI ( P11ENI )
     ,.P04ENI ( P04ENI ) ,.P12ENI ( P12ENI ) ,.P20ENI ( P20ENI ) ,.P05ENI ( P05ENI )
     ,.P13ENI ( P13ENI ) ,.P21ENI ( P21ENI ) ,.P06ENI ( P06ENI ) ,.P14ENI ( P14ENI )
     ,.P22ENI ( P22ENI ) ,.P30ENI ( P30ENI ) ,.P00DIN ( P00DIN ) ,.P01DIN ( P01DIN )
     ,.P02DIN ( P02DIN ) ,.P10DIN ( P10DIN ) ,.P03DIN ( P03DIN ) ,.P11DIN ( P11DIN )
     ,.P04DIN ( P04DIN ) ,.P12DIN ( P12DIN ) ,.P20DIN ( P20DIN ) ,.P05DIN ( P05DIN )
     ,.P13DIN ( P13DIN ) ,.P21DIN ( P21DIN ) ,.P06DIN ( P06DIN ) ,.P14DIN ( P14DIN )
     ,.P22DIN ( P22DIN ) ,.P30DIN ( P30DIN ) ,.P01SELIN ( P01SELIN ) ,.P03SELIN ( P03SELIN )
     ,.P11SELIN ( P11SELIN ) ,.P04SELIN ( P04SELIN ) ,.P15ENO ( P15ENO )
     ,.P23ENO ( P23ENO ) ,.P31ENO ( P31ENO ) ,.P16ENO ( P16ENO ) ,.P24ENO ( P24ENO )
     ,.P40ENO ( P40ENO ) ,.P17ENO ( P17ENO ) ,.P25ENO ( P25ENO ) ,.P41ENO ( P41ENO )
     ,.P15DOUT ( P15DOUT ) ,.P23DOUT ( P23DOUT ) ,.P31DOUT ( P31DOUT )
     ,.P16DOUT ( P16DOUT ) ,.P24DOUT ( P24DOUT ) ,.P40DOUT ( P40DOUT )
     ,.P17DOUT ( P17DOUT ) ,.P25DOUT ( P25DOUT ) ,.P41DOUT ( P41DOUT )
     ,.P15ENI ( P15ENI ) ,.P23ENI ( P23ENI ) ,.P31ENI ( P31ENI ) ,.P16ENI ( P16ENI )
     ,.P24ENI ( P24ENI ) ,.P40ENI ( P40ENI ) ,.P17ENI ( P17ENI ) ,.P25ENI ( P25ENI )
     ,.P41ENI ( P41ENI ) ,.P15DIN ( P15DIN ) ,.P23DIN ( P23DIN ) ,.P31DIN ( P31DIN )
     ,.P16DIN ( P16DIN ) ,.P24DIN ( P24DIN ) ,.P40DIN ( P40DIN ) ,.P17DIN ( P17DIN )
     ,.P25DIN ( P25DIN ) ,.P41DIN ( P41DIN ) ,.P10SELIN ( P10SELIN ) ,.P13SELIN ( P13SELIN )
     ,.P14SELIN ( P14SELIN ) ,.P15SELIN ( P15SELIN ) ,.P16SELIN ( P16SELIN )
     ,.P17SELIN ( P17SELIN ) ,.P26ENO ( P26ENO ) ,.P42ENO ( P42ENO ) ,.P50ENO ( P50ENO )
     ,.P27ENO ( P27ENO ) ,.P43ENO ( P43ENO ) ,.P51ENO ( P51ENO ) ,.P26DOUT ( P26DOUT )
     ,.P42DOUT ( P42DOUT ) ,.P50DOUT ( P50DOUT ) ,.P27DOUT ( P27DOUT )
     ,.P43DOUT ( P43DOUT ) ,.P51DOUT ( P51DOUT ) ,.P26ENI ( P26ENI ) ,.P42ENI ( P42ENI )
     ,.P50ENI ( P50ENI ) ,.P27ENI ( P27ENI ) ,.P43ENI ( P43ENI ) ,.P51ENI ( P51ENI )
     ,.P26DIN ( P26DIN ) ,.P42DIN ( P42DIN ) ,.P50DIN ( P50DIN ) ,.P27DIN ( P27DIN )
     ,.P43DIN ( P43DIN ) ,.P51DIN ( P51DIN ) ,.P52ENO ( P52ENO ) ,.P60ENO ( P60ENO )
     ,.P53ENO ( P53ENO ) ,.P61ENO ( P61ENO ) ,.DGEN07 ( DGEN07 ) ,.P54ENO ( P54ENO )
     ,.P62ENO ( P62ENO ) ,.P70ENO ( P70ENO ) ,.P55ENO ( P55ENO ) ,.P63ENO ( P63ENO )
     ,.P71ENO ( P71ENO ) ,.P52DOUT ( P52DOUT ) ,.P60DOUT ( P60DOUT ) ,.P53DOUT ( P53DOUT )
     ,.P61DOUT ( P61DOUT ) ,.P54DOUT ( P54DOUT ) ,.P62DOUT ( P62DOUT )
     ,.P70DOUT ( P70DOUT ) ,.P55DOUT ( P55DOUT ) ,.P63DOUT ( P63DOUT )
     ,.P71DOUT ( P71DOUT ) ,.P52ENI ( P52ENI ) ,.P60ENI ( P60ENI ) ,.P53ENI ( P53ENI )
     ,.P61ENI ( P61ENI ) ,.DGEN01 ( DGEN01 ) ,.P54ENI ( P54ENI ) ,.P62ENI ( P62ENI )
     ,.P70ENI ( P70ENI ) ,.P55ENI ( P55ENI ) ,.P63ENI ( P63ENI ) ,.P71ENI ( P71ENI )
     ,.P52DIN ( P52DIN ) ,.P60DIN ( P60DIN ) ,.P53DIN ( P53DIN ) ,.P61DIN ( P61DIN )
     ,.P54DIN ( P54DIN ) ,.P62DIN ( P62DIN ) ,.P70DIN ( P70DIN ) ,.DGEN00 ( DGEN00 )
     ,.P55DIN ( P55DIN ) ,.P63DIN ( P63DIN ) ,.P71DIN ( P71DIN ) ,.P55SELIN ( P55SELIN )
     ,.P72ENO ( P72ENO ) ,.P73ENO ( P73ENO ) ,.P74ENO ( P74ENO ) ,.P75ENO ( P75ENO )
     ,.P76ENO ( P76ENO ) ,.AD_DB3 ( AD_DB3 ) ,.P77ENO ( P77ENO ) ,.P72DOUT ( P72DOUT )
     ,.P73DOUT ( P73DOUT ) ,.P74DOUT ( P74DOUT ) ,.P75DOUT ( P75DOUT )
     ,.P76DOUT ( P76DOUT ) ,.P77DOUT ( P77DOUT ) ,.P72ENI ( P72ENI ) ,.P73ENI ( P73ENI )
     ,.P74ENI ( P74ENI ) ,.P75ENI ( P75ENI ) ,.P76ENI ( P76ENI ) ,.P77ENI ( P77ENI )
     ,.AD_DB5 ( AD_DB5 ) ,.P72DIN ( P72DIN ) ,.P73DIN ( P73DIN ) ,.P74DIN ( P74DIN )
     ,.ADRD_B ( ADRD_B ) ,.P75DIN ( P75DIN ) ,.P76DIN ( P76DIN ) ,.P77DIN ( P77DIN )
     ,.ADSH_B ( ADSH_B ) ,.P120ENO ( P120ENO ) ,.P120DOUT ( P120DOUT )
     ,.P120ENI ( P120ENI ) ,.P120DIN ( P120DIN ) ,.P130ENO ( P130ENO )
     ,.P130DOUT ( P130DOUT ) ,.P137ENI ( P137ENI ) ,.P137DIN ( P137DIN )
     ,.P140ENO ( P140ENO ) ,.P141ENO ( P141ENO ) ,.P146ENO ( P146ENO )
     ,.P147ENO ( P147ENO ) ,.P140DOUT ( P140DOUT ) ,.P141DOUT ( P141DOUT )
     ,.P146DOUT ( P146DOUT ) ,.P147DOUT ( P147DOUT ) ,.P140ENI ( P140ENI )
     ,.P141ENI ( P141ENI ) ,.P146ENI ( P146ENI ) ,.P147ENI ( P147ENI )
     ,.P140DIN ( P140DIN ) ,.P141DIN ( P141DIN ) ,.P146DIN ( P146DIN )
     ,.P147DIN ( P147DIN ) ,.P00PUON ( P00PUON ) ,.P01PUON ( P01PUON )
     ,.P02PUON ( P02PUON ) ,.P10PUON ( P10PUON ) ,.P03PUON ( P03PUON )
     ,.P11PUON ( P11PUON ) ,.P04PUON ( P04PUON ) ,.P12PUON ( P12PUON )
     ,.P05PUON ( P05PUON ) ,.P13PUON ( P13PUON ) ,.ADINT_B ( ADINT_B )
     ,.P06PUON ( P06PUON ) ,.P14PUON ( P14PUON ) ,.P30PUON ( P30PUON )
     ,.P15PUON ( P15PUON ) ,.P31PUON ( P31PUON ) ,.P16PUON ( P16PUON )
     ,.P40PUON ( P40PUON ) ,.P17PUON ( P17PUON ) ,.P41PUON ( P41PUON )
     ,.P42PUON ( P42PUON ) ,.P50PUON ( P50PUON ) ,.P43PUON ( P43PUON )
     ,.P51PUON ( P51PUON ) ,.P52PUON ( P52PUON ) ,.P53PUON ( P53PUON )
     ,.P54PUON ( P54PUON ) ,.P70PUON ( P70PUON ) ,.P55PUON ( P55PUON )
     ,.P71PUON ( P71PUON ) ,.P72PUON ( P72PUON ) ,.P75PUON ( P75PUON )
     ,.P76PUON ( P76PUON ) ,.P77PUON ( P77PUON ) ,.P120PUON ( P120PUON )
     ,.P140PUON ( P140PUON ) ,.P141PUON ( P141PUON ) ,.P146PUON ( P146PUON )
     ,.P147PUON ( P147PUON ) ,.PIO00 ( PIO00 ) ,.PIO01 ( PIO01 ) ,.PIO02 ( PIO02 )
     ,.PIO10 ( PIO10 ) ,.PIO03 ( PIO03 ) ,.PIO11 ( PIO11 ) ,.PIO04 ( PIO04 )
     ,.PIO12 ( PIO12 ) ,.PIO20 ( PIO20 ) ,.PIO05 ( PIO05 ) ,.PIO13 ( PIO13 )
     ,.PIO21 ( PIO21 ) ,.PIO06 ( PIO06 ) ,.PIO14 ( PIO14 ) ,.PIO22 ( PIO22 )
     ,.PIO30 ( PIO30 ) ,.PIO15 ( PIO15 ) ,.PIO23 ( PIO23 ) ,.PIO31 ( PIO31 )
     ,.PIO16 ( PIO16 ) ,.PIO24 ( PIO24 ) ,.PIO40 ( PIO40 ) ,.PIO17 ( PIO17 )
     ,.PIO25 ( PIO25 ) ,.PIO41 ( PIO41 ) ,.PIO26 ( PIO26 ) ,.PIO42 ( PIO42 )
     ,.PIO50 ( PIO50 ) ,.PIO27 ( PIO27 ) ,.PIO43 ( PIO43 ) ,.PIO51 ( PIO51 )
     ,.PIO52 ( PIO52 ) ,.PIO60 ( PIO60 ) ,.PIO53 ( PIO53 ) ,.PIO61 ( PIO61 )
     ,.PIO54 ( PIO54 ) ,.PIO62 ( PIO62 ) ,.PIO70 ( PIO70 ) ,.PIO55 ( PIO55 )
     ,.PIO63 ( PIO63 ) ,.PIO71 ( PIO71 ) ,.PIO72 ( PIO72 ) ,.PIO73 ( PIO73 )
     ,.PIO74 ( PIO74 ) ,.PIO75 ( PIO75 ) ,.PIO76 ( PIO76 ) ,.PIO77 ( PIO77 )
     ,.PIO120 ( PIO120 ) ,.PIO121 ( PIO121 ) ,.PIO122 ( PIO122 ) ,.PIO130 ( PIO130 )
     ,.PIO123 ( PIO123 ) ,.PIO124 ( PIO124 ) ,.PIO140 ( PIO140 ) ,.PIO137 ( PIO137 )
     ,.PIO141 ( PIO141 ) ,.PIO146 ( PIO146 ) ,.PIO147 ( PIO147 ) ,.PSEUDOANI09 ( PSEUDOANI09 )
     ,.PSEUDOANI17 ( PSEUDOANI17 ) ,.PSEUDOANI08 ( PSEUDOANI08 ) ,.PSEUDOANI16 ( PSEUDOANI16 )
     ,.PSEUDOANI07 ( PSEUDOANI07 ) ,.PSEUDOANI15 ( PSEUDOANI15 ) ,.PSEUDOANI06 ( PSEUDOANI06 )
     ,.PSEUDOANI14 ( PSEUDOANI14 ) ,.PSEUDOANI05 ( PSEUDOANI05 ) ,.PSEUDOANI13 ( PSEUDOANI13 )
     ,.PSEUDOANI04 ( PSEUDOANI04 ) ,.PSEUDOANI12 ( PSEUDOANI12 ) ,.PSEUDOANI03 ( PSEUDOANI03 )
     ,.PSEUDOANI11 ( PSEUDOANI11 ) ,.PSEUDOANI02 ( PSEUDOANI02 ) ,.PSEUDOANI10 ( PSEUDOANI10 )
     ,.PSEUDOANI01 ( PSEUDOANI01 ) ,.PSEUDOANI00 ( PSEUDOANI00 ) ,.PSEUDOANI19 ( PSEUDOANI19 )
     ,.PSEUDOANI18 ( PSEUDOANI18 ) ,.AD_DB9 ( AD_DB9 ) ,.AD_DB8 ( AD_DB8 )
     ,.AD_DB7 ( AD_DB7 ) ,.AD_DB6 ( AD_DB6 ) ,.AD_DB4 ( AD_DB4 ) ,.AD_DB2 ( AD_DB2 )
     ,.AD_DB1 ( AD_DB1 ) ,.AD_DB0 ( AD_DB0 ) ,.ADCS_B ( ADCS_B ) ,.AD_A4 ( AD_A4 )
     ,.AD_A3 ( AD_A3 ) ,.AD_A2 ( AD_A2 ) ,.AD_A1 ( AD_A1 ) ,.AD_A0 ( AD_A0 )
     ,.ADGSELMOD ( ADGSELMOD ) ,.ADVSELMOD0_I ( ADVSELMOD0_I ) ,.ADVSELMOD1_I ( ADVSELMOD1_I )
     ,.DGEN06 ( DGEN06 ) ,.DGEN05 ( DGEN05 ) ,.DGEN04 ( DGEN04 ) ,.DGEN03 ( DGEN03 )
     ,.DGEN02 ( DGEN02 )
  ) ;
  // Refer to /home/product/div-micom-ice/data/proj/78K0R/Common/ICEMacro/tags/SS3rd_V1_0_32/ice_top_SS3rd.v
  ICE_TOP ice (
    .CLK30MHZ_GB ( CLK30MHZ_GB ) ,.A19 ( A19 ) ,.A18 ( A18 ) ,.A17 ( A17 )
     ,.A16 ( A16 ) ,.A15 ( A15 ) ,.A14 ( A14 ) ,.A13 ( A13 ) ,.A12 ( A12 )
     ,.A11 ( A11 ) ,.A10 ( A10 ) ,.A9 ( A9 ) ,.A8 ( A8 ) ,.A7 ( A7 ) ,.A6 ( A6 )
     ,.A5 ( A5 ) ,.A4 ( A4 ) ,.A3 ( A3 ) ,.A2 ( A2 ) ,.DW37 ( DW37 ) ,.DW29 ( DW29 )
     ,.PA13 ( PA13 ) ,.DW36 ( DW36 ) ,.DW28 ( DW28 ) ,.PA12 ( PA12 ) ,.DW35 ( DW35 )
     ,.DW27 ( DW27 ) ,.DW19 ( DW19 ) ,.PA11 ( PA11 ) ,.DW34 ( DW34 ) ,.DW26 ( DW26 )
     ,.DW18 ( DW18 ) ,.PA10 ( PA10 ) ,.DW33 ( DW33 ) ,.DW25 ( DW25 ) ,.DW17 ( DW17 )
     ,.DDIS ( DDIS ) ,.DW32 ( DW32 ) ,.DW24 ( DW24 ) ,.DW16 ( DW16 ) ,.DW31 ( DW31 )
     ,.DW23 ( DW23 ) ,.DW15 ( DW15 ) ,.DW30 ( DW30 ) ,.DW22 ( DW22 ) ,.DW14 ( DW14 )
     ,.DW21 ( DW21 ) ,.DW13 ( DW13 ) ,.ALT1 ( ALT1 ) ,.DW20 ( DW20 ) ,.DW12 ( DW12 )
     ,.DW11 ( DW11 ) ,.DW10 ( DW10 ) ,.DW9 ( DW9 ) ,.PA5 ( PA5 ) ,.PC1 ( PC1 )
     ,.DW8 ( DW8 ) ,.PA4 ( PA4 ) ,.PC0 ( PC0 ) ,.DW7 ( DW7 ) ,.DIS ( DIS )
     ,.PA3 ( PA3 ) ,.DW6 ( DW6 ) ,.PA2 ( PA2 ) ,.DW5 ( DW5 ) ,.DW4 ( DW4 )
     ,.DW3 ( DW3 ) ,.DW2 ( DW2 ) ,.DW1 ( DW1 ) ,.MA9 ( MA9 ) ,.DW0 ( DW0 )
     ,.MA8 ( MA8 ) ,.BEU2 ( BEU2 ) ,.MA12 ( MA12 ) ,.BEU1 ( BEU1 ) ,.MA11 ( MA11 )
     ,.BEU0 ( BEU0 ) ,.MA10 ( MA10 ) ,.READ ( READ ) ,.MRG00 ( MRG00 )
     ,.MRG01 ( MRG01 ) ,.MRG10 ( MRG10 ) ,.MRG11 ( MRG11 ) ,.MRG12 ( MRG12 )
     ,.WWR ( WWR ) ,.CLKSEL1 ( CLKSEL1 ) ,.RDCLKP1 ( RDCLKP1 ) ,.FCLK ( FCLK1 )
     ,.PA19 ( PA19 ) ,.PC11 ( PC11 ) ,.PROGI ( PROGI ) ,.USBA1 ( USBA1 )
     ,.CER ( CER ) ,.MA2 ( MA2 ) ,.SER ( SER ) ,.CE0 ( CE0 ) ,.AF6 ( AF6 )
     ,.DA4 ( DA4 ) ,.CE1 ( CE1 ) ,.AF7 ( AF7 ) ,.DA5 ( DA5 ) ,.EXA ( EXA )
     ,.WED ( WED ) ,.EXCH ( EXCH ) ,.MDW0 ( MDW0 ) ,.FLMD0 ( pull_down1 )
     ,.SELRO1 ( SELRO1 ) ,.BRSAM ( BRSAM ) ,.ICEWAITMEM ( ICEWAITMEM )
     ,.ICENOECC ( ICENOECC ) ,.ICEFLERR ( ICEFLERR ) ,.RO137 ( RO137 )
     ,.RO129 ( RO129 ) ,.EXMA3 ( EXMA3 ) ,.RO136 ( RO136 ) ,.RO128 ( RO128 )
     ,.EXMA2 ( EXMA2 ) ,.RO135 ( RO135 ) ,.RO127 ( RO127 ) ,.RO119 ( RO119 )
     ,.EXMA1 ( EXMA1 ) ,.RO134 ( RO134 ) ,.RO126 ( RO126 ) ,.RO118 ( RO118 )
     ,.EXMA0 ( EXMA0 ) ,.RO133 ( RO133 ) ,.RO125 ( RO125 ) ,.RO117 ( RO117 )
     ,.RO037 ( RO037 ) ,.RO029 ( RO029 ) ,.RO132 ( RO132 ) ,.RO124 ( RO124 )
     ,.RO116 ( RO116 ) ,.RO036 ( RO036 ) ,.RO028 ( RO028 ) ,.RO131 ( RO131 )
     ,.RO123 ( RO123 ) ,.RO115 ( RO115 ) ,.RO035 ( RO035 ) ,.RO027 ( RO027 )
     ,.RO019 ( RO019 ) ,.RO130 ( RO130 ) ,.RO122 ( RO122 ) ,.RO114 ( RO114 )
     ,.RO034 ( RO034 ) ,.RO026 ( RO026 ) ,.RO018 ( RO018 ) ,.RO121 ( RO121 )
     ,.RO113 ( RO113 ) ,.RO033 ( RO033 ) ,.RO025 ( RO025 ) ,.RO017 ( RO017 )
     ,.RO120 ( RO120 ) ,.RO112 ( RO112 ) ,.RO032 ( RO032 ) ,.RO024 ( RO024 )
     ,.RO016 ( RO016 ) ,.RO111 ( RO111 ) ,.RO031 ( RO031 ) ,.RO023 ( RO023 )
     ,.RO015 ( RO015 ) ,.RO110 ( RO110 ) ,.RO030 ( RO030 ) ,.RO022 ( RO022 )
     ,.RO014 ( RO014 ) ,.RO19 ( RO19 ) ,.RO18 ( RO18 ) ,.RO17 ( RO17 )
     ,.RO09 ( RO09 ) ,.RO16 ( RO16 ) ,.RO08 ( RO08 ) ,.RO15 ( RO15 ) ,.RO07 ( RO07 )
     ,.RO14 ( RO14 ) ,.RO06 ( RO06 ) ,.RO13 ( RO13 ) ,.RO05 ( RO05 ) ,.RO12 ( RO12 )
     ,.RO04 ( RO04 ) ,.RO11 ( RO11 ) ,.RO03 ( RO03 ) ,.MDW9 ( MDW9 ) ,.RO10 ( RO10 )
     ,.RO02 ( RO02 ) ,.MDW8 ( MDW8 ) ,.RO021 ( RO021 ) ,.RO013 ( RO013 )
     ,.RO020 ( RO020 ) ,.RO012 ( RO012 ) ,.CPURD ( CPURD ) ,.RO011 ( RO011 )
     ,.RO010 ( RO010 ) ,.RO01 ( RO01 ) ,.MDW7 ( MDW7 ) ,.RO00 ( RO00 )
     ,.MDW6 ( MDW6 ) ,.WAITFL2 ( WAITFL2 ) ,.SLFLASH ( SLFLASH ) ,.TMEMA14 ( TMEMA14 )
     ,.GDRAMWR ( GDRAMWR ) ,.CIBPID31 ( CIBPID31 ) ,.CIBPID23 ( CIBPID23 )
     ,.CIBPID15 ( CIBPID15 ) ,.CIBPID30 ( CIBPID30 ) ,.CIBPID22 ( CIBPID22 )
     ,.CIBPID14 ( CIBPID14 ) ,.CIBPID29 ( CIBPID29 ) ,.CIBPID28 ( CIBPID28 )
     ,.CIBPID27 ( CIBPID27 ) ,.CIBPID19 ( CIBPID19 ) ,.CIBPID26 ( CIBPID26 )
     ,.CIBPID18 ( CIBPID18 ) ,.CIBPID25 ( CIBPID25 ) ,.CIBPID17 ( CIBPID17 )
     ,.CIBPID24 ( CIBPID24 ) ,.CIBPID16 ( CIBPID16 ) ,.CIBPID21 ( CIBPID21 )
     ,.CIBPID13 ( CIBPID13 ) ,.CIBPID20 ( CIBPID20 ) ,.CIBPID12 ( CIBPID12 )
     ,.CIBPID11 ( CIBPID11 ) ,.CIBPID10 ( CIBPID10 ) ,.CIBPID9 ( CIBPID9 )
     ,.CIBPID8 ( CIBPID8 ) ,.CIBPID7 ( CIBPID7 ) ,.CIBPID6 ( CIBPID6 )
     ,.CIBPID5 ( CIBPID5 ) ,.CIBPID4 ( CIBPID4 ) ,.CIBPID3 ( CIBPID3 )
     ,.CIBPID2 ( CIBPID2 ) ,.CIBPID1 ( CIBPID1 ) ,.CIBPID0 ( CIBPID0 )
     ,.CPUPID31 ( CPUPID31 ) ,.CPUPID23 ( CPUPID23 ) ,.CPUPID15 ( CPUPID15 )
     ,.CPUPID30 ( CPUPID30 ) ,.CPUPID22 ( CPUPID22 ) ,.CPUPID14 ( CPUPID14 )
     ,.CPUPID29 ( CPUPID29 ) ,.CPUPID28 ( CPUPID28 ) ,.CPUPID27 ( CPUPID27 )
     ,.CPUPID19 ( CPUPID19 ) ,.CPUPID26 ( CPUPID26 ) ,.CPUPID18 ( CPUPID18 )
     ,.CPUPID25 ( CPUPID25 ) ,.CPUPID17 ( CPUPID17 ) ,.CPUPID24 ( CPUPID24 )
     ,.CPUPID16 ( CPUPID16 ) ,.CPUPID21 ( CPUPID21 ) ,.CPUPID13 ( CPUPID13 )
     ,.CPUPID20 ( CPUPID20 ) ,.CPUPID12 ( CPUPID12 ) ,.CPUPID11 ( CPUPID11 )
     ,.CPUPID10 ( CPUPID10 ) ,.CPUPID9 ( CPUPID9 ) ,.CPUPID8 ( CPUPID8 )
     ,.CPUPID7 ( CPUPID7 ) ,.CPUPID6 ( CPUPID6 ) ,.CPUPID5 ( CPUPID5 )
     ,.CPUPID4 ( CPUPID4 ) ,.CPUPID3 ( CPUPID3 ) ,.CPUPID2 ( CPUPID2 )
     ,.CPUPID1 ( CPUPID1 ) ,.CPUMASK ( CPUMASK ) ,.CPUPID0 ( CPUPID0 )
     ,.ICEIFA31 ( ICEIFA31 ) ,.ICEIFA23 ( ICEIFA23 ) ,.ICEIFA15 ( ICEIFA15 )
     ,.ICEIFA30 ( ICEIFA30 ) ,.ICEIFA22 ( ICEIFA22 ) ,.ICEIFA14 ( ICEIFA14 )
     ,.ICEIFA29 ( ICEIFA29 ) ,.ICEIFA28 ( ICEIFA28 ) ,.ICEIFA27 ( ICEIFA27 )
     ,.ICEIFA19 ( ICEIFA19 ) ,.ICEIFA26 ( ICEIFA26 ) ,.ICEIFA18 ( ICEIFA18 )
     ,.ICEIFA25 ( ICEIFA25 ) ,.ICEIFA17 ( ICEIFA17 ) ,.ICEIFA24 ( ICEIFA24 )
     ,.ICEIFA16 ( ICEIFA16 ) ,.ICEIFA21 ( ICEIFA21 ) ,.ICEIFA13 ( ICEIFA13 )
     ,.ICEDOA29 ( ICEDO29 ) ,.ICEIFA20 ( ICEIFA20 ) ,.ICEIFA12 ( ICEIFA12 )
     ,.ICEDOA28 ( ICEDO28 ) ,.ICEIFA11 ( ICEIFA11 ) ,.ICEDOA27 ( ICEDO27 )
     ,.ICEDOA19 ( ICEDO19 ) ,.ICEIFA10 ( ICEIFA10 ) ,.ICEDOA26 ( ICEDO26 )
     ,.ICEDOA18 ( ICEDO18 ) ,.ICEIFA9 ( ICEIFA9 ) ,.ICEIFA8 ( ICEIFA8 )
     ,.ICEIFA7 ( ICEIFA7 ) ,.ICEIFA6 ( ICEIFA6 ) ,.ICEIFA5 ( ICEIFA5 )
     ,.ICEDOA9 ( ICEDO9 ) ,.ICEIFA4 ( ICEIFA4 ) ,.ICEDOA8 ( ICEDO8 ) ,.ICEIFA3 ( ICEIFA3 )
     ,.ICEDOA7 ( ICEDO7 ) ,.ICEIFA2 ( ICEIFA2 ) ,.ICEDOA6 ( ICEDO6 ) ,.ICEIFA1 ( ICEIFA1 )
     ,.ICEDOA5 ( ICEDO5 ) ,.ICEIFA0 ( ICEIFA0 ) ,.ICEDOA4 ( ICEDO4 ) ,.ICEDI31 ( ICEDI31 )
     ,.ICEDI23 ( ICEDI23 ) ,.ICEDI15 ( ICEDI15 ) ,.IDADR11 ( IDADR11 )
     ,.ICEDI30 ( ICEDI30 ) ,.ICEDI22 ( ICEDI22 ) ,.ICEDI14 ( ICEDI14 )
     ,.IDADR10 ( IDADR10 ) ,.ICEDI29 ( ICEDI29 ) ,.IDADR25 ( IDADR25 )
     ,.IDADR17 ( IDADR17 ) ,.ICEDI28 ( ICEDI28 ) ,.IDADR24 ( IDADR24 )
     ,.IDADR16 ( IDADR16 ) ,.ICEDI27 ( ICEDI27 ) ,.ICEDI19 ( ICEDI19 )
     ,.IDADR31 ( IDADR31 ) ,.IDADR23 ( IDADR23 ) ,.IDADR15 ( IDADR15 )
     ,.ICEDI26 ( ICEDI26 ) ,.ICEDI18 ( ICEDI18 ) ,.IDADR30 ( IDADR30 )
     ,.IDADR22 ( IDADR22 ) ,.IDADR14 ( IDADR14 ) ,.ICEDI25 ( ICEDI25 )
     ,.ICEDI17 ( ICEDI17 ) ,.IDADR21 ( IDADR21 ) ,.IDADR13 ( IDADR13 )
     ,.ICEDI24 ( ICEDI24 ) ,.ICEDI16 ( ICEDI16 ) ,.IDADR20 ( IDADR20 )
     ,.IDADR12 ( IDADR12 ) ,.ICEDI21 ( ICEDI21 ) ,.ICEDI13 ( ICEDI13 )
     ,.ICEDI20 ( ICEDI20 ) ,.ICEDI12 ( ICEDI12 ) ,.ICEDI11 ( ICEDI11 )
     ,.ICEDI10 ( ICEDI10 ) ,.ICEDI9 ( ICEDI9 ) ,.IDADR7 ( IDADR7 ) ,.ICEDI8 ( ICEDI8 )
     ,.IDADR6 ( IDADR6 ) ,.ICEDI7 ( ICEDI7 ) ,.IDADR5 ( IDADR5 ) ,.ICEDI6 ( ICEDI6 )
     ,.IDADR4 ( IDADR4 ) ,.ICEDI5 ( ICEDI5 ) ,.IDADR3 ( IDADR3 ) ,.ICEDI4 ( ICEDI4 )
     ,.IDADR2 ( IDADR2 ) ,.ICEDI3 ( ICEDI3 ) ,.IDADR1 ( IDADR1 ) ,.ICEDI2 ( ICEDI2 )
     ,.IDADR0 ( IDADR0 ) ,.ICEDI1 ( ICEDI1 ) ,.ICEDI0 ( ICEDI0 ) ,.ICEWR ( ICEWR )
     ,.ICEDOP31 ( ICEDOP31 ) ,.ICEDOP23 ( ICEDOP23 ) ,.ICEDOP15 ( ICEDOP15 )
     ,.ICEDOP30 ( ICEDOP30 ) ,.ICEDOP22 ( ICEDOP22 ) ,.ICEDOP14 ( ICEDOP14 )
     ,.ICEDOP29 ( ICEDOP29 ) ,.ICEDOP28 ( ICEDOP28 ) ,.ICEDOP27 ( ICEDOP27 )
     ,.ICEDOP19 ( ICEDOP19 ) ,.ICEDOP26 ( ICEDOP26 ) ,.ICEDOP18 ( ICEDOP18 )
     ,.ICEDOP25 ( ICEDOP25 ) ,.ICEDOP17 ( ICEDOP17 ) ,.ICEDOP24 ( ICEDOP24 )
     ,.ICEDOP16 ( ICEDOP16 ) ,.ICEDOP21 ( ICEDOP21 ) ,.ICEDOP13 ( ICEDOP13 )
     ,.ICEDOP20 ( ICEDOP20 ) ,.ICEDOP12 ( ICEDOP12 ) ,.ICEDOP11 ( ICEDOP11 )
     ,.ICEDOP10 ( ICEDOP10 ) ,.ICEDOP9 ( ICEDOP9 ) ,.ICEDOP8 ( ICEDOP8 )
     ,.ICEDOP7 ( ICEDOP7 ) ,.ICEDOP6 ( ICEDOP6 ) ,.ICEDOP5 ( ICEDOP5 )
     ,.ICEDOP4 ( ICEDOP4 ) ,.ICEDOP3 ( ICEDOP3 ) ,.ICEDOP2 ( ICEDOP2 )
     ,.ICEDOP1 ( ICEDOP1 ) ,.ICEDOP0 ( ICEDOP0 ) ,.ICEDOA31 ( ICEDO31 )
     ,.ICEDOA23 ( ICEDO23 ) ,.ICEDOA15 ( ICEDO15 ) ,.ICEDOA30 ( ICEDO30 )
     ,.ICEDOA22 ( ICEDO22 ) ,.ICEDOA14 ( ICEDO14 ) ,.ICEDOA25 ( ICEDO25 )
     ,.ICEDOA17 ( ICEDO17 ) ,.ICEDOA24 ( ICEDO24 ) ,.ICEDOA16 ( ICEDO16 )
     ,.ICEDOA21 ( ICEDO21 ) ,.ICEDOA13 ( ICEDO13 ) ,.ICEDOA20 ( ICEDO20 )
     ,.ICEDOA12 ( ICEDO12 ) ,.ICEDOA11 ( ICEDO11 ) ,.ICEDOA10 ( ICEDO10 )
     ,.ICEDOA3 ( ICEDO3 ) ,.ICEDOA2 ( ICEDO2 ) ,.ICEDOA1 ( ICEDO1 ) ,.ICEDOA0 ( ICEDO0 )
     ,.VDDLEV7 ( VDDLEV7 ) ,.VDDLEV6 ( VDDLEV6 ) ,.VDDLEV5 ( VDDLEV5 )
     ,.VDDLEV4 ( VDDLEV4 ) ,.VDDLEV3 ( VDDLEV3 ) ,.VDDLEV2 ( VDDLEV2 )
     ,.VDDLEV1 ( VDDLEV1 ) ,.VDDLEV0 ( VDDLEV0 ) ,.USBIFWR ( USBIFWR )
     ,.ICECSGREGU ( ICECSGREGU ) ,.POCRESB ( POCRESB ) ,.TARRESB ( RESINB )
     ,.CPUPRCLK2 ( pull_down3 ) ,.CPUTMCLK ( CPUTMCLK ) ,.CPUTSCLK ( CPUTSCLK )
     ,.CPURCLK1SEL ( pull_down2 ) ,.CLK60MHZ ( CLK60MHZ ) ,.CLK60MHZLOCK ( CLK60MHZLOCK )
     ,.CPUMCLK ( CPUMCLK ) ,.CPUSCLK ( CPUSCLK ) ,.CPURCLK1 ( CPURCLK1 )
     ,.CPURCLK2 ( CPURCLK2 ) ,.CPURCLK3 ( CPURCLK3 ) ,.SOFTBRK ( SBANDOCD )
     ,.SVINTACK ( SVINTACK ) ,.STBRELESV ( STBRELESV ) ,.SVI ( SVI ) ,.SVMODI ( SVMODI )
     ,.SVMODIPERI1 ( SVMODIPERI1 ) ,.SVMODIPERI2 ( SVMODIPERI2 ) ,.SVVCOUT7 ( SVVCOUT7 )
     ,.SVVCOUT6 ( SVVCOUT6 ) ,.SVVCOUT5 ( SVVCOUT5 ) ,.SVVCOUT4 ( SVVCOUT4 )
     ,.SVVCOUT3 ( SVVCOUT3 ) ,.SVVCOUT2 ( SVVCOUT2 ) ,.SVVCOUT1 ( SVVCOUT1 )
     ,.SVVCOUT0 ( SVVCOUT0 ) ,.SVMODOPBRK ( SVMODOPBRK ) ,.IDADR29 ( IDADR29 )
     ,.IDADR28 ( IDADR28 ) ,.IDADR27 ( IDADR27 ) ,.IDADR19 ( IDADR19 )
     ,.IDADR26 ( IDADR26 ) ,.IDADR18 ( IDADR18 ) ,.IDADR9 ( IDADR9 ) ,.IDADR8 ( IDADR8 )
     ,.PERISVIB ( PERISVIB ) ,.FLSIZE3 ( FLSIZE3 ) ,.FLSIZE2 ( FLSIZE2 )
     ,.FLSIZE1 ( FLSIZE1 ) ,.FLSIZE0 ( FLSIZE0 ) ,.RAMSIZE7 ( RAMSIZE7 )
     ,.RAMSIZE6 ( RAMSIZE6 ) ,.RAMSIZE5 ( RAMSIZE5 ) ,.RAMSIZE4 ( RAMSIZE4 )
     ,.RAMSIZE3 ( RAMSIZE3 ) ,.RAMSIZE2 ( RAMSIZE2 ) ,.RAMSIZE1 ( RAMSIZE1 )
     ,.RAMSIZE0 ( RAMSIZE0 ) ,.BFSIZE3 ( BFSIZE3 ) ,.BFSIZE2 ( BFSIZE2 )
     ,.BFSIZE1 ( BFSIZE1 ) ,.BFSIZE0 ( BFSIZE0 ) ,.BMSIZE3 ( BMSIZE3 )
     ,.BMSIZE2 ( BMSIZE2 ) ,.BMSIZE1 ( BMSIZE1 ) ,.BMSIZE0 ( BMSIZE0 )
     ,.DFSIZE1 ( DFSIZE1 ) ,.DFSIZE0 ( DFSIZE0 ) ,.PSEUDOON31 ( PSEUDOON31 )
     ,.PSEUDOON23 ( PSEUDOON23 ) ,.PSEUDOON15 ( PSEUDOON15 ) ,.PSEUDOON30 ( PSEUDOON30 )
     ,.PSEUDOON22 ( PSEUDOON22 ) ,.PSEUDOON14 ( PSEUDOON14 ) ,.PSEUDOON29 ( PSEUDOON29 )
     ,.PSEUDOON28 ( PSEUDOON28 ) ,.PSEUDOON27 ( PSEUDOON27 ) ,.PSEUDOON19 ( PSEUDOON19 )
     ,.PSEUDOON26 ( PSEUDOON26 ) ,.PSEUDOON18 ( PSEUDOON18 ) ,.PSEUDOON25 ( PSEUDOON25 )
     ,.PSEUDOON17 ( PSEUDOON17 ) ,.PSEUDOON24 ( PSEUDOON24 ) ,.PSEUDOON16 ( PSEUDOON16 )
     ,.PSEUDOON21 ( PSEUDOON21 ) ,.PSEUDOON13 ( PSEUDOON13 ) ,.PSEUDOON20 ( PSEUDOON20 )
     ,.PSEUDOON12 ( PSEUDOON12 ) ,.PSEUDOON11 ( PSEUDOON11 ) ,.PSEUDOON10 ( PSEUDOON10 )
     ,.PSEUDOON9 ( PSEUDOON9 ) ,.PSEUDOON8 ( PSEUDOON8 ) ,.PSEUDOON7 ( PSEUDOON7 )
     ,.PSEUDOON6 ( PSEUDOON6 ) ,.PSEUDOON5 ( PSEUDOON5 ) ,.PSEUDOON4 ( PSEUDOON4 )
     ,.PSEUDOON3 ( PSEUDOON3 ) ,.PSEUDOON2 ( PSEUDOON2 ) ,.PSEUDOON1 ( PSEUDOON1 )
     ,.PSEUDOON0 ( PSEUDOON0 ) ,.PSEUDOANI09 ( PSEUDOANI09 ) ,.PSEUDOANI17 ( PSEUDOANI17 )
     ,.PSEUDOANI08 ( PSEUDOANI08 ) ,.PSEUDOANI16 ( PSEUDOANI16 ) ,.PSEUDOANI07 ( PSEUDOANI07 )
     ,.PSEUDOANI15 ( PSEUDOANI15 ) ,.PSEUDOANI06 ( PSEUDOANI06 ) ,.PSEUDOANI14 ( PSEUDOANI14 )
     ,.PSEUDOANI05 ( PSEUDOANI05 ) ,.PSEUDOANI13 ( PSEUDOANI13 ) ,.PSEUDOANI04 ( PSEUDOANI04 )
     ,.PSEUDOANI12 ( PSEUDOANI12 ) ,.PSEUDOANI03 ( PSEUDOANI03 ) ,.PSEUDOANI11 ( PSEUDOANI11 )
     ,.PSEUDOANI02 ( PSEUDOANI02 ) ,.PSEUDOANI10 ( PSEUDOANI10 ) ,.PSEUDOANI01 ( PSEUDOANI01 )
     ,.PSEUDOANI00 ( PSEUDOANI00 ) ,.PSEUDOANI19 ( PSEUDOANI19 ) ,.PSEUDOANI18 ( PSEUDOANI18 )
     ,.ICEMSKDBG ( ICEMSKDBG ) ,.ICEMSKWAIT ( ICEMSKWAIT ) ,.ICEMSKNMI ( ICEMSKNMI )
     ,.ICEMSKTRAP ( ICEMSKTRAP ) ,.ICEMSKWDT ( ICEMKWDT ) ,.ICEMSKLVI ( ICEMKLVI )
     ,.ICEMSKRETRY ( ICEMSKRETRY ) ,.MDR_RAM15 ( MDRRAM15 ) ,.MDR_RAM14 ( MDRRAM14 )
     ,.MDR_RAM13 ( MDRRAM13 ) ,.MDR_RAM12 ( MDRRAM12 ) ,.MDR_RAM11 ( MDRRAM11 )
     ,.MDR_RAM10 ( MDRRAM10 ) ,.MDR_RAM9 ( MDRRAM9 ) ,.MDR_RAM8 ( MDRRAM8 )
     ,.MDR_RAM7 ( MDRRAM7 ) ,.MDR_RAM6 ( MDRRAM6 ) ,.MDR_RAM5 ( MDRRAM5 )
     ,.MDR_RAM4 ( MDRRAM4 ) ,.MDR_RAM3 ( MDRRAM3 ) ,.MDR_RAM2 ( MDRRAM2 )
     ,.MDR_RAM1 ( MDRRAM1 ) ,.MDR_RAM0 ( MDRRAM0 ) ,.CPUWR ( CPUWR ) ,.WDOP ( WDOP )
     ,.SVMOD ( SVMOD ) ,.SVMODF ( SVMODF ) ,.STAGEADR1 ( STAGEADR1 ) ,.STAGEADR0 ( STAGEADR0 )
     ,.PCWAITF ( PCWAITF ) ,.SKIPEXE ( SKIPEXE ) ,.FCHRAM ( FCHRAM ) ,.FLREAD ( FLREAD )
     ,.IMDR10 ( IMDR10 ) ,.FLREADB3 ( FLREADB3 ) ,.FLREADB2 ( FLREADB2 )
     ,.FLREADB1 ( FLREADB1 ) ,.FLREADB0 ( FLREADB0 ) ,.CPURSOUTB ( RESETB )
     ,.BASECK ( FCLK_ICE ) ,.PREFIX ( PREFIX ) ,.WAITEXM ( pull_down0 )
     ,.OCDWAIT ( OCDWAIT ) ,.BRAMEN ( pull_up0 ) ,.BFA ( BFA ) ,.BFAEN ( pull_up1 )
     ,.INTACK ( INTACK ) ,.DMAACK ( DMAACK ) ,.SLEXM ( SLEXM ) ,.IDPOP ( IDPOP )
     ,.MDW10 ( MDW10 ) ,.IMDR2 ( IMDR2 ) ,.SPINC ( SPINC ) ,.SPDEC ( SPDEC )
     ,.SPREL ( SPREL ) ,.CPUMISAL ( CPUMISAL ) ,.SLMEM ( SLMEM ) ,.FLSPMD ( FLSPM )
     ,.STPST ( STPST ) ,.HLTST ( HLTST ) ,.MA15 ( MA15 ) ,.MA14 ( MA14 )
     ,.MA13 ( MA13 ) ,.MA7 ( MA7 ) ,.MA6 ( MA6 ) ,.MA5 ( MA5 ) ,.MA4 ( MA4 )
     ,.MA3 ( MA3 ) ,.MA1 ( MA1 ) ,.MA0 ( MA0 ) ,.MDW15 ( MDW15 ) ,.IMDR7 ( IMDR7 )
     ,.MDW14 ( MDW14 ) ,.IMDR6 ( IMDR6 ) ,.MDW13 ( MDW13 ) ,.IMDR5 ( IMDR5 )
     ,.MDW12 ( MDW12 ) ,.IMDR4 ( IMDR4 ) ,.MDW11 ( MDW11 ) ,.IMDR3 ( IMDR3 )
     ,.MDW5 ( MDW5 ) ,.MDW4 ( MDW4 ) ,.MDW3 ( MDW3 ) ,.MDW2 ( MDW2 ) ,.MDW1 ( MDW1 )
     ,.PA18 ( PA18 ) ,.PC10 ( PC10 ) ,.PA17 ( PA17 ) ,.PA16 ( PA16 ) ,.PA15 ( PA15 )
     ,.PA14 ( PA14 ) ,.PA9 ( PA9 ) ,.PC5 ( PC5 ) ,.PA8 ( PA8 ) ,.PC4 ( PC4 )
     ,.PA7 ( PA7 ) ,.PC3 ( PC3 ) ,.PA6 ( PA6 ) ,.PC2 ( PC2 ) ,.PC19 ( PC19 )
     ,.PC18 ( PC18 ) ,.PC17 ( PC17 ) ,.PC16 ( PC16 ) ,.PC15 ( PC15 ) ,.PC14 ( PC14 )
     ,.PC13 ( PC13 ) ,.PC12 ( PC12 ) ,.PC9 ( PC9 ) ,.PC8 ( PC8 ) ,.PC7 ( PC7 )
     ,.PC6 ( PC6 ) ,.IMDR15 ( IMDR15 ) ,.IMDR14 ( IMDR14 ) ,.IMDR13 ( IMDR13 )
     ,.IMDR12 ( IMDR12 ) ,.IMDR11 ( IMDR11 ) ,.IMDR9 ( IMDR9 ) ,.IMDR8 ( IMDR8 )
     ,.IMDR1 ( IMDR1 ) ,.IMDR0 ( IMDR0 ) ,.SLBMEM ( SLBMEM ) ,.SYSRSOUTB ( SYSRSOUTB )
     ,.PONRESB ( PONRESB ) ,.CPUPRCLK3 ( CPUPRCLK3 ) ,.LOCKFAIL5 ( LOCK64FAIL )
     ,.LOCKFAIL6 ( LOCK48FAIL ) ,.LOCKFAIL7 ( LOCKHROSCFAIL ) ,.LOCKFAIL8 ( pull_down7 )
     ,.LOCKFAIL9 ( pull_down8 ) ,.LOCKFAIL10 ( pull_down9 ) ,.LOCKFAIL11 ( pull_down10 )
     ,.LOCKFAIL12 ( pull_down11 ) ,.LOCKFAIL20 ( pull_down19 ) ,.LOCKFAIL13 ( pull_down12 )
     ,.LOCKFAIL21 ( pull_down20 ) ,.LOCKFAIL14 ( pull_down13 ) ,.LOCKFAIL22 ( pull_down21 )
     ,.LOCKFAIL30 ( pull_down29 ) ,.LOCKFAIL15 ( pull_down14 ) ,.LOCKFAIL23 ( pull_down22 )
     ,.LOCKFAIL16 ( pull_down15 ) ,.LOCKFAIL24 ( pull_down23 ) ,.LOCKFAIL17 ( pull_down16 )
     ,.LOCKFAIL25 ( pull_down24 ) ,.LOCKFAIL18 ( pull_down17 ) ,.LOCKFAIL26 ( pull_down25 )
     ,.LOCKFAIL19 ( pull_down18 ) ,.LOCKFAIL27 ( pull_down26 ) ,.LOCKFAIL28 ( pull_down27 )
     ,.LOCKFAIL29 ( pull_down28 ) ,.IDVER31 ( IDVER31 ) ,.IDVER23 ( IDVER23 )
     ,.IDVER15 ( IDVER15 ) ,.IDVER30 ( IDVER30 ) ,.IDVER22 ( IDVER22 )
     ,.IDVER14 ( IDVER14 ) ,.IDVER29 ( IDVER29 ) ,.IDVER28 ( IDVER28 )
     ,.IDVER27 ( IDVER27 ) ,.IDVER19 ( IDVER19 ) ,.IDVER26 ( IDVER26 )
     ,.IDVER18 ( IDVER18 ) ,.IDVER25 ( IDVER25 ) ,.IDVER17 ( IDVER17 )
     ,.IDVER24 ( IDVER24 ) ,.IDVER16 ( IDVER16 ) ,.IDVER21 ( IDVER21 )
     ,.IDVER13 ( IDVER13 ) ,.IDVER20 ( IDVER20 ) ,.IDVER12 ( IDVER12 )
     ,.IDVER11 ( IDVER11 ) ,.IDVER10 ( IDVER10 ) ,.IDVER9 ( IDVER9 ) ,.IDVER8 ( IDVER8 )
     ,.IDVER7 ( IDVER7 ) ,.IDVER6 ( IDVER6 ) ,.IDVER5 ( IDVER5 ) ,.IDVER4 ( IDVER4 )
     ,.IDVER3 ( IDVER3 ) ,.IDVER2 ( IDVER2 ) ,.IDVER1 ( IDVER1 ) ,.IDVER0 ( IDVER0 )
     ,.ADDRTD144 ( ADDRTD144 ) ,.ADDRTD136 ( ADDRTD136 ) ,.ADDRTD128 ( ADDRTD128 )
     ,.ADDRTD143 ( ADDRTD143 ) ,.ADDRTD135 ( ADDRTD135 ) ,.ADDRTD127 ( ADDRTD127 )
     ,.ADDRTD119 ( ADDRTD119 ) ,.ADDRTD142 ( ADDRTD142 ) ,.ADDRTD134 ( ADDRTD134 )
     ,.ADDRTD126 ( ADDRTD126 ) ,.ADDRTD118 ( ADDRTD118 ) ,.ADDRTD141 ( ADDRTD141 )
     ,.ADDRTD133 ( ADDRTD133 ) ,.ADDRTD125 ( ADDRTD125 ) ,.ADDRTD117 ( ADDRTD117 )
     ,.ADDRTD109 ( ADDRTD109 ) ,.ADDRTD140 ( ADDRTD140 ) ,.ADDRTD132 ( ADDRTD132 )
     ,.ADDRTD124 ( ADDRTD124 ) ,.ADDRTD116 ( ADDRTD116 ) ,.ADDRTD108 ( ADDRTD108 )
     ,.ADDRTD139 ( ADDRTD139 ) ,.ADDRTD138 ( ADDRTD138 ) ,.ADDRTD137 ( ADDRTD137 )
     ,.ADDRTD129 ( ADDRTD129 ) ,.ADDRTD131 ( ADDRTD131 ) ,.ADDRTD123 ( ADDRTD123 )
     ,.ADDRTD115 ( ADDRTD115 ) ,.ADDRTD107 ( ADDRTD107 ) ,.ADDRTD130 ( ADDRTD130 )
     ,.ADDRTD122 ( ADDRTD122 ) ,.ADDRTD114 ( ADDRTD114 ) ,.ADDRTD106 ( ADDRTD106 )
     ,.ADDRTD121 ( ADDRTD121 ) ,.ADDRTD113 ( ADDRTD113 ) ,.ADDRTD105 ( ADDRTD105 )
     ,.ADDRTD120 ( ADDRTD120 ) ,.ADDRTD112 ( ADDRTD112 ) ,.ADDRTD104 ( ADDRTD104 )
     ,.ADDRTD111 ( ADDRTD111 ) ,.ADDRTD103 ( ADDRTD103 ) ,.ADDRTD110 ( ADDRTD110 )
     ,.ADDRTD102 ( ADDRTD102 ) ,.ADDRTD101 ( ADDRTD101 ) ,.ADDRTD100 ( ADDRTD100 )
     ,.ADDRTD99 ( ADDRTD99 ) ,.ADDRTD98 ( ADDRTD98 ) ,.ADDRTD97 ( ADDRTD97 )
     ,.ADDRTD89 ( ADDRTD89 ) ,.ADDRTD96 ( ADDRTD96 ) ,.ADDRTD88 ( ADDRTD88 )
     ,.ADDRTD95 ( ADDRTD95 ) ,.ADDRTD87 ( ADDRTD87 ) ,.ADDRTD79 ( ADDRTD79 )
     ,.ADDRTD94 ( ADDRTD94 ) ,.ADDRTD86 ( ADDRTD86 ) ,.ADDRTD78 ( ADDRTD78 )
     ,.ADDRTD93 ( ADDRTD93 ) ,.ADDRTD85 ( ADDRTD85 ) ,.ADDRTD77 ( ADDRTD77 )
     ,.ADDRTD69 ( ADDRTD69 ) ,.ADDRTD92 ( ADDRTD92 ) ,.ADDRTD84 ( ADDRTD84 )
     ,.ADDRTD76 ( ADDRTD76 ) ,.ADDRTD68 ( ADDRTD68 ) ,.ADDRTD91 ( ADDRTD91 )
     ,.ADDRTD83 ( ADDRTD83 ) ,.ADDRTD75 ( ADDRTD75 ) ,.ADDRTD67 ( ADDRTD67 )
     ,.ADDRTD59 ( ADDRTD59 ) ,.ADDRTD90 ( ADDRTD90 ) ,.ADDRTD82 ( ADDRTD82 )
     ,.ADDRTD74 ( ADDRTD74 ) ,.ADDRTD66 ( ADDRTD66 ) ,.ADDRTD58 ( ADDRTD58 )
     ,.ADDRTD81 ( ADDRTD81 ) ,.ADDRTD73 ( ADDRTD73 ) ,.ADDRTD65 ( ADDRTD65 )
     ,.ADDRTD57 ( ADDRTD57 ) ,.ADDRTD49 ( ADDRTD49 ) ,.ADDRTD80 ( ADDRTD80 )
     ,.ADDRTD72 ( ADDRTD72 ) ,.ADDRTD64 ( ADDRTD64 ) ,.ADDRTD56 ( ADDRTD56 )
     ,.ADDRTD48 ( ADDRTD48 ) ,.ADDRTD71 ( ADDRTD71 ) ,.ADDRTD63 ( ADDRTD63 )
     ,.ADDRTD55 ( ADDRTD55 ) ,.ADDRTD47 ( ADDRTD47 ) ,.ADDRTD39 ( ADDRTD39 )
     ,.ADDRTD70 ( ADDRTD70 ) ,.ADDRTD62 ( ADDRTD62 ) ,.ADDRTD54 ( ADDRTD54 )
     ,.ADDRTD46 ( ADDRTD46 ) ,.ADDRTD38 ( ADDRTD38 ) ,.ADDRTD61 ( ADDRTD61 )
     ,.ADDRTD53 ( ADDRTD53 ) ,.ADDRTD45 ( ADDRTD45 ) ,.ADDRTD37 ( ADDRTD37 )
     ,.ADDRTD29 ( ADDRTD29 ) ,.ADDRTD60 ( ADDRTD60 ) ,.ADDRTD52 ( ADDRTD52 )
     ,.ADDRTD44 ( ADDRTD44 ) ,.ADDRTD36 ( ADDRTD36 ) ,.ADDRTD28 ( ADDRTD28 )
     ,.ADDRTD51 ( ADDRTD51 ) ,.ADDRTD43 ( ADDRTD43 ) ,.ADDRTD35 ( ADDRTD35 )
     ,.ADDRTD27 ( ADDRTD27 ) ,.ADDRTD19 ( ADDRTD19 ) ,.ADDRTD50 ( ADDRTD50 )
     ,.ADDRTD42 ( ADDRTD42 ) ,.ADDRTD34 ( ADDRTD34 ) ,.ADDRTD26 ( ADDRTD26 )
     ,.ADDRTD18 ( ADDRTD18 ) ,.ADDRTD41 ( ADDRTD41 ) ,.ADDRTD33 ( ADDRTD33 )
     ,.ADDRTD25 ( ADDRTD25 ) ,.ADDRTD17 ( ADDRTD17 ) ,.ADDRTD40 ( ADDRTD40 )
     ,.ADDRTD32 ( ADDRTD32 ) ,.ADDRTD24 ( ADDRTD24 ) ,.ADDRTD16 ( ADDRTD16 )
     ,.ADDRTD31 ( ADDRTD31 ) ,.ADDRTD23 ( ADDRTD23 ) ,.ADDRTD15 ( ADDRTD15 )
     ,.ADDRTD30 ( ADDRTD30 ) ,.ADDRTD22 ( ADDRTD22 ) ,.ADDRTD14 ( ADDRTD14 )
     ,.ADDRTD21 ( ADDRTD21 ) ,.ADDRTD13 ( ADDRTD13 ) ,.ADDRTD20 ( ADDRTD20 )
     ,.ADDRTD12 ( ADDRTD12 ) ,.ADDRTD11 ( ADDRTD11 ) ,.ADDRTD10 ( ADDRTD10 )
     ,.ADDRTD9 ( ADDRTD9 ) ,.ADDRTD8 ( ADDRTD8 ) ,.ADDRTD7 ( ADDRTD7 )
     ,.ADDRTD6 ( ADDRTD6 ) ,.ADDRTD5 ( ADDRTD5 ) ,.ADDRTD4 ( ADDRTD4 )
     ,.ADDRTD3 ( ADDRTD3 ) ,.ADDRTD2 ( ADDRTD2 ) ,.ADDRTD1 ( ADDRTD1 )
     ,.ADDRPINRD ( ADDRPINRD ) ,.ADDRPINMD ( ADDRPINMD ) ,.ADDRPINLV ( ADDRPINLV )
     ,.TP144D3 ( pull_down172 ) ,.TP136D3 ( pull_down204 ) ,.TP128D3 ( pull_down236 )
     ,.TP144D2 ( pull_down173 ) ,.TP136D2 ( pull_down205 ) ,.TP128D2 ( pull_down237 )
     ,.TP144D1 ( pull_down174 ) ,.TP136D1 ( pull_down206 ) ,.TP128D1 ( pull_down238 )
     ,.TP144D0 ( pull_down175 ) ,.TP136D0 ( pull_down207 ) ,.TP128D0 ( pull_down239 )
     ,.TP143D3 ( pull_down176 ) ,.TP135D3 ( pull_down208 ) ,.TP127D3 ( pull_down240 )
     ,.TP119D3 ( pull_down272 ) ,.TP143D2 ( pull_down177 ) ,.TP135D2 ( pull_down209 )
     ,.TP127D2 ( pull_down241 ) ,.TP119D2 ( pull_down273 ) ,.TP143D1 ( pull_down178 )
     ,.TP135D1 ( pull_down210 ) ,.TP127D1 ( pull_down242 ) ,.TP119D1 ( pull_down274 )
     ,.TP143D0 ( pull_down179 ) ,.TP135D0 ( pull_down211 ) ,.TP127D0 ( pull_down243 )
     ,.TP119D0 ( pull_down275 ) ,.TP142D3 ( pull_down180 ) ,.TP134D3 ( pull_down212 )
     ,.TP126D3 ( pull_down244 ) ,.TP118D3 ( pull_down276 ) ,.TP142D2 ( pull_down181 )
     ,.TP134D2 ( pull_down213 ) ,.TP126D2 ( pull_down245 ) ,.TP118D2 ( pull_down277 )
     ,.TP142D1 ( pull_down182 ) ,.TP134D1 ( pull_down214 ) ,.TP126D1 ( pull_down246 )
     ,.TP118D1 ( pull_down278 ) ,.TP142D0 ( pull_down183 ) ,.TP134D0 ( pull_down215 )
     ,.TP126D0 ( pull_down247 ) ,.TP118D0 ( pull_down279 ) ,.TP141D3 ( pull_down184 )
     ,.TP133D3 ( pull_down216 ) ,.TP125D3 ( pull_down248 ) ,.TP117D3 ( pull_down280 )
     ,.TP109D3 ( pull_down312 ) ,.TP141D2 ( pull_down185 ) ,.TP133D2 ( pull_down217 )
     ,.TP125D2 ( pull_down249 ) ,.TP117D2 ( pull_down281 ) ,.TP109D2 ( pull_down313 )
     ,.TP141D1 ( pull_down186 ) ,.TP133D1 ( pull_down218 ) ,.TP125D1 ( pull_down250 )
     ,.TP117D1 ( pull_down282 ) ,.TP109D1 ( pull_down314 ) ,.TP141D0 ( pull_down187 )
     ,.TP133D0 ( pull_down219 ) ,.TP125D0 ( pull_down251 ) ,.TP117D0 ( pull_down283 )
     ,.TP109D0 ( pull_down315 ) ,.TP140D3 ( pull_down188 ) ,.TP132D3 ( pull_down220 )
     ,.TP124D3 ( pull_down252 ) ,.TP116D3 ( pull_down284 ) ,.TP108D3 ( pull_down316 )
     ,.TP140D2 ( pull_down189 ) ,.TP132D2 ( pull_down221 ) ,.TP124D2 ( pull_down253 )
     ,.TP116D2 ( pull_down285 ) ,.TP108D2 ( pull_down317 ) ,.TP140D1 ( pull_down190 )
     ,.TP132D1 ( pull_down222 ) ,.TP124D1 ( pull_down254 ) ,.TP116D1 ( pull_down286 )
     ,.TP108D1 ( pull_down318 ) ,.TP140D0 ( pull_down191 ) ,.TP132D0 ( pull_down223 )
     ,.TP124D0 ( pull_down255 ) ,.TP116D0 ( pull_down287 ) ,.TP108D0 ( pull_down319 )
     ,.TP139D3 ( pull_down192 ) ,.TP139D2 ( pull_down193 ) ,.TP139D1 ( pull_down194 )
     ,.TP139D0 ( pull_down195 ) ,.TP138D3 ( pull_down196 ) ,.TP138D2 ( pull_down197 )
     ,.TP138D1 ( pull_down198 ) ,.TP138D0 ( pull_down199 ) ,.TP137D3 ( pull_down200 )
     ,.TP129D3 ( pull_down232 ) ,.TP137D2 ( pull_down201 ) ,.TP129D2 ( pull_down233 )
     ,.TP137D1 ( pull_down202 ) ,.TP129D1 ( pull_down234 ) ,.TP137D0 ( pull_down203 )
     ,.TP129D0 ( pull_down235 ) ,.TP131D3 ( pull_down224 ) ,.TP123D3 ( pull_down256 )
     ,.TP115D3 ( pull_down288 ) ,.TP107D3 ( pull_down320 ) ,.TP131D2 ( pull_down225 )
     ,.TP123D2 ( pull_down257 ) ,.TP115D2 ( pull_down289 ) ,.TP107D2 ( pull_down321 )
     ,.TP131D1 ( pull_down226 ) ,.TP123D1 ( pull_down258 ) ,.TP115D1 ( pull_down290 )
     ,.TP107D1 ( pull_down322 ) ,.TP131D0 ( pull_down227 ) ,.TP123D0 ( pull_down259 )
     ,.TP115D0 ( pull_down291 ) ,.TP107D0 ( pull_down323 ) ,.TP130D3 ( pull_down228 )
     ,.TP122D3 ( pull_down260 ) ,.TP114D3 ( pull_down292 ) ,.TP106D3 ( pull_down324 )
     ,.TP130D2 ( pull_down229 ) ,.TP122D2 ( pull_down261 ) ,.TP114D2 ( pull_down293 )
     ,.TP106D2 ( pull_down325 ) ,.TP130D1 ( pull_down230 ) ,.TP122D1 ( pull_down262 )
     ,.TP114D1 ( pull_down294 ) ,.TP106D1 ( pull_down326 ) ,.TP130D0 ( pull_down231 )
     ,.TP122D0 ( pull_down263 ) ,.TP114D0 ( pull_down295 ) ,.TP106D0 ( pull_down327 )
     ,.TP121D3 ( pull_down264 ) ,.TP113D3 ( pull_down296 ) ,.TP105D3 ( pull_down328 )
     ,.TP121D2 ( pull_down265 ) ,.TP113D2 ( pull_down297 ) ,.TP105D2 ( pull_down329 )
     ,.TP121D1 ( pull_down266 ) ,.TP113D1 ( pull_down298 ) ,.TP105D1 ( pull_down330 )
     ,.TP121D0 ( pull_down267 ) ,.TP113D0 ( pull_down299 ) ,.TP105D0 ( pull_down331 )
     ,.TP120D3 ( pull_down268 ) ,.TP112D3 ( pull_down300 ) ,.TP104D3 ( pull_down332 )
     ,.TP120D2 ( pull_down269 ) ,.TP112D2 ( pull_down301 ) ,.TP104D2 ( pull_down333 )
     ,.EROMWRB ( EROMWRB ) ,.TP120D1 ( pull_down270 ) ,.TP112D1 ( pull_down302 )
     ,.TP104D1 ( pull_down334 ) ,.TP120D0 ( pull_down271 ) ,.TP112D0 ( pull_down303 )
     ,.TP104D0 ( pull_down335 ) ,.TP111D3 ( pull_down304 ) ,.TP103D3 ( pull_down336 )
     ,.TP111D2 ( pull_down305 ) ,.TP103D2 ( pull_down337 ) ,.TP111D1 ( pull_down306 )
     ,.TP103D1 ( pull_down338 ) ,.TP111D0 ( pull_down307 ) ,.TP103D0 ( pull_down339 )
     ,.TP110D3 ( pull_down308 ) ,.TP102D3 ( pull_down340 ) ,.TP110D2 ( pull_down309 )
     ,.TP102D2 ( pull_down341 ) ,.TP110D1 ( pull_down310 ) ,.TP102D1 ( pull_down342 )
     ,.TP110D0 ( pull_down311 ) ,.TP102D0 ( pull_down343 ) ,.TP101D3 ( pull_down344 )
     ,.TP101D2 ( pull_down345 ) ,.TP101D1 ( pull_down346 ) ,.TP101D0 ( pull_down347 )
     ,.TP100D3 ( pull_down348 ) ,.TP100D2 ( pull_down349 ) ,.TP100D1 ( pull_down350 )
     ,.TP100D0 ( pull_down351 ) ,.TP99D3 ( pull_down352 ) ,.TP99D2 ( pull_down353 )
     ,.TP99D1 ( pull_down354 ) ,.TP99D0 ( pull_down355 ) ,.TP98D3 ( pull_down356 )
     ,.TP98D2 ( pull_down357 ) ,.TP98D1 ( pull_down358 ) ,.TP98D0 ( pull_down359 )
     ,.TP97D3 ( pull_down360 ) ,.TP89D3 ( pull_down392 ) ,.TP97D2 ( pull_down361 )
     ,.TP89D2 ( pull_down393 ) ,.TP97D1 ( pull_down362 ) ,.TP89D1 ( pull_down394 )
     ,.TP97D0 ( pull_down363 ) ,.TP89D0 ( pull_down395 ) ,.TP96D3 ( pull_down364 )
     ,.TP88D3 ( pull_down396 ) ,.TP96D2 ( pull_down365 ) ,.TP88D2 ( pull_down397 )
     ,.TP96D1 ( pull_down366 ) ,.TP88D1 ( pull_down398 ) ,.TP96D0 ( pull_down367 )
     ,.TP88D0 ( pull_down399 ) ,.TP95D3 ( pull_down368 ) ,.TP87D3 ( pull_down400 )
     ,.TP79D3 ( pull_down432 ) ,.TP95D2 ( pull_down369 ) ,.TP87D2 ( pull_down401 )
     ,.TP79D2 ( pull_down433 ) ,.TP95D1 ( pull_down370 ) ,.TP87D1 ( pull_down402 )
     ,.TP79D1 ( pull_down434 ) ,.TP95D0 ( pull_down371 ) ,.TP87D0 ( pull_down403 )
     ,.TP79D0 ( pull_down435 ) ,.TP94D3 ( pull_down372 ) ,.TP86D3 ( pull_down404 )
     ,.TP78D3 ( pull_down436 ) ,.TP94D2 ( pull_down373 ) ,.TP86D2 ( pull_down405 )
     ,.TP78D2 ( pull_down437 ) ,.TP94D1 ( pull_down374 ) ,.TP86D1 ( pull_down406 )
     ,.TP78D1 ( pull_down438 ) ,.TP94D0 ( pull_down375 ) ,.TP86D0 ( pull_down407 )
     ,.TP78D0 ( pull_down439 ) ,.TP93D3 ( pull_down376 ) ,.TP85D3 ( pull_down408 )
     ,.TP77D3 ( pull_down440 ) ,.TP69D3 ( pull_down472 ) ,.TP93D2 ( pull_down377 )
     ,.TP85D2 ( pull_down409 ) ,.TP77D2 ( pull_down441 ) ,.TP69D2 ( pull_down473 )
     ,.TP93D1 ( pull_down378 ) ,.TP85D1 ( pull_down410 ) ,.TP77D1 ( pull_down442 )
     ,.TP69D1 ( pull_down474 ) ,.TP93D0 ( pull_down379 ) ,.TP85D0 ( pull_down411 )
     ,.TP77D0 ( pull_down443 ) ,.TP69D0 ( pull_down475 ) ,.TP92D3 ( pull_down380 )
     ,.TP84D3 ( pull_down412 ) ,.TP76D3 ( pull_down444 ) ,.TP68D3 ( pull_down476 )
     ,.TP92D2 ( pull_down381 ) ,.TP84D2 ( pull_down413 ) ,.TP76D2 ( pull_down445 )
     ,.TP68D2 ( pull_down477 ) ,.TP92D1 ( pull_down382 ) ,.TP84D1 ( pull_down414 )
     ,.TP76D1 ( pull_down446 ) ,.TP68D1 ( pull_down478 ) ,.TP92D0 ( pull_down383 )
     ,.TP84D0 ( pull_down415 ) ,.TP76D0 ( pull_down447 ) ,.TP68D0 ( pull_down479 )
     ,.TP91D3 ( pull_down384 ) ,.TP83D3 ( pull_down416 ) ,.TP75D3 ( pull_down448 )
     ,.TP67D3 ( pull_down480 ) ,.TP59D3 ( pull_down512 ) ,.TP91D2 ( pull_down385 )
     ,.TP83D2 ( pull_down417 ) ,.TP75D2 ( pull_down449 ) ,.TP67D2 ( pull_down481 )
     ,.TP59D2 ( pull_down513 ) ,.TP91D1 ( pull_down386 ) ,.TP83D1 ( pull_down418 )
     ,.TP75D1 ( pull_down450 ) ,.TP67D1 ( pull_down482 ) ,.TP59D1 ( pull_down514 )
     ,.TP91D0 ( pull_down387 ) ,.TP83D0 ( pull_down419 ) ,.TP75D0 ( pull_down451 )
     ,.TP67D0 ( pull_down483 ) ,.TP59D0 ( pull_down515 ) ,.TP90D3 ( pull_down388 )
     ,.TP82D3 ( pull_down420 ) ,.TP74D3 ( pull_down452 ) ,.TP66D3 ( pull_down484 )
     ,.TP58D3 ( pull_down516 ) ,.TP90D2 ( pull_down389 ) ,.TP82D2 ( pull_down421 )
     ,.TP74D2 ( pull_down453 ) ,.TP66D2 ( pull_down485 ) ,.TP58D2 ( pull_down517 )
     ,.TP90D1 ( pull_down390 ) ,.TP82D1 ( pull_down422 ) ,.TP74D1 ( pull_down454 )
     ,.TP66D1 ( pull_down486 ) ,.TP58D1 ( pull_down518 ) ,.TP90D0 ( pull_down391 )
     ,.TP82D0 ( pull_down423 ) ,.TP74D0 ( pull_down455 ) ,.TP66D0 ( pull_down487 )
     ,.TP58D0 ( pull_down519 ) ,.TP81D3 ( pull_down424 ) ,.TP73D3 ( pull_down456 )
     ,.TP65D3 ( pull_down488 ) ,.TP57D3 ( pull_down520 ) ,.TP49D3 ( pull_down552 )
     ,.TP81D2 ( pull_down425 ) ,.TP73D2 ( pull_down457 ) ,.TP65D2 ( pull_down489 )
     ,.TP57D2 ( pull_down521 ) ,.TP49D2 ( pull_down553 ) ,.TP81D1 ( pull_down426 )
     ,.TP73D1 ( pull_down458 ) ,.TP65D1 ( pull_down490 ) ,.TP57D1 ( pull_down522 )
     ,.TP49D1 ( pull_down554 ) ,.TP81D0 ( pull_down427 ) ,.TP73D0 ( pull_down459 )
     ,.TP65D0 ( pull_down491 ) ,.TP57D0 ( pull_down523 ) ,.TP49D0 ( pull_down555 )
     ,.TP80D3 ( pull_down428 ) ,.TP72D3 ( pull_down460 ) ,.TP64D3 ( pull_down492 )
     ,.TP56D3 ( pull_down524 ) ,.TP48D3 ( pull_down556 ) ,.TP80D2 ( pull_down429 )
     ,.TP72D2 ( pull_down461 ) ,.TP64D2 ( pull_down493 ) ,.TP56D2 ( pull_down525 )
     ,.TP48D2 ( pull_down557 ) ,.TP80D1 ( pull_down430 ) ,.TP72D1 ( pull_down462 )
     ,.TP64D1 ( pull_down494 ) ,.TP56D1 ( pull_down526 ) ,.TP48D1 ( pull_down558 )
     ,.TP80D0 ( pull_down431 ) ,.TP72D0 ( pull_down463 ) ,.TP64D0 ( pull_down495 )
     ,.TP56D0 ( pull_down527 ) ,.TP48D0 ( pull_down559 ) ,.TP71D3 ( pull_down464 )
     ,.TP63D3 ( pull_down496 ) ,.TP55D3 ( pull_down528 ) ,.TP47D3 ( pull_down560 )
     ,.TP39D3 ( pull_down592 ) ,.TP71D2 ( pull_down465 ) ,.TP63D2 ( pull_down497 )
     ,.TP55D2 ( pull_down529 ) ,.TP47D2 ( pull_down561 ) ,.TP39D2 ( pull_down593 )
     ,.TP71D1 ( pull_down466 ) ,.TP63D1 ( pull_down498 ) ,.TP55D1 ( pull_down530 )
     ,.TP47D1 ( pull_down562 ) ,.TP39D1 ( pull_down594 ) ,.TP71D0 ( pull_down467 )
     ,.TP63D0 ( pull_down499 ) ,.TP55D0 ( pull_down531 ) ,.TP47D0 ( pull_down563 )
     ,.TP39D0 ( pull_down595 ) ,.TP70D3 ( pull_down468 ) ,.TP62D3 ( pull_down500 )
     ,.TP54D3 ( pull_down532 ) ,.TP46D3 ( pull_down564 ) ,.TP38D3 ( pull_down596 )
     ,.TP70D2 ( pull_down469 ) ,.TP62D2 ( pull_down501 ) ,.TP54D2 ( pull_down533 )
     ,.TP46D2 ( pull_down565 ) ,.TP38D2 ( pull_down597 ) ,.TP70D1 ( pull_down470 )
     ,.TP62D1 ( pull_down502 ) ,.TP54D1 ( pull_down534 ) ,.TP46D1 ( pull_down566 )
     ,.TP38D1 ( pull_down598 ) ,.TP70D0 ( pull_down471 ) ,.TP62D0 ( pull_down503 )
     ,.TP54D0 ( pull_down535 ) ,.TP46D0 ( pull_down567 ) ,.TP38D0 ( pull_down599 )
     ,.TP61D3 ( pull_down504 ) ,.TP53D3 ( pull_down536 ) ,.TP45D3 ( pull_down568 )
     ,.TP37D3 ( pull_down600 ) ,.TP29D3 ( pull_down632 ) ,.TP61D2 ( pull_down505 )
     ,.TP53D2 ( pull_down537 ) ,.TP45D2 ( pull_down569 ) ,.TP37D2 ( pull_down601 )
     ,.TP29D2 ( pull_down633 ) ,.TP61D1 ( pull_down506 ) ,.TP53D1 ( pull_down538 )
     ,.TP45D1 ( pull_down570 ) ,.TP37D1 ( pull_down602 ) ,.TP29D1 ( pull_down634 )
     ,.TP61D0 ( pull_down507 ) ,.TP53D0 ( pull_down539 ) ,.TP45D0 ( pull_down571 )
     ,.TP37D0 ( pull_down603 ) ,.TP29D0 ( pull_down635 ) ,.TP60D3 ( pull_down508 )
     ,.TP52D3 ( pull_down540 ) ,.TP44D3 ( pull_down572 ) ,.TP36D3 ( pull_down604 )
     ,.TP28D3 ( pull_down636 ) ,.TP60D2 ( pull_down509 ) ,.TP52D2 ( pull_down541 )
     ,.TP44D2 ( pull_down573 ) ,.TP36D2 ( pull_down605 ) ,.TP28D2 ( pull_down637 )
     ,.TP60D1 ( pull_down510 ) ,.TP52D1 ( pull_down542 ) ,.TP44D1 ( pull_down574 )
     ,.TP36D1 ( pull_down606 ) ,.TP28D1 ( pull_down638 ) ,.TP60D0 ( pull_down511 )
     ,.TP52D0 ( pull_down543 ) ,.TP44D0 ( pull_down575 ) ,.TP36D0 ( pull_down607 )
     ,.TP28D0 ( pull_down639 ) ,.TP51D3 ( pull_down544 ) ,.TP43D3 ( pull_down576 )
     ,.TP35D3 ( pull_down608 ) ,.TP27D3 ( pull_down640 ) ,.TP19D3 ( pull_down672 )
     ,.TP51D2 ( pull_down545 ) ,.TP43D2 ( pull_down577 ) ,.TP35D2 ( pull_down609 )
     ,.TP27D2 ( pull_down641 ) ,.TP19D2 ( pull_down673 ) ,.TP51D1 ( pull_down546 )
     ,.TP43D1 ( pull_down578 ) ,.TP35D1 ( pull_down610 ) ,.TP27D1 ( pull_down642 )
     ,.TP19D1 ( pull_down674 ) ,.TP51D0 ( pull_down547 ) ,.TP43D0 ( pull_down579 )
     ,.TP35D0 ( pull_down611 ) ,.TP27D0 ( pull_down643 ) ,.TP19D0 ( pull_down675 )
     ,.TP50D3 ( pull_down548 ) ,.TP42D3 ( pull_down580 ) ,.TP34D3 ( pull_down612 )
     ,.TP26D3 ( pull_down644 ) ,.TP18D3 ( pull_down676 ) ,.TP50D2 ( pull_down549 )
     ,.TP42D2 ( pull_down581 ) ,.TP34D2 ( pull_down613 ) ,.TP26D2 ( pull_down645 )
     ,.TP18D2 ( pull_down677 ) ,.TP50D1 ( pull_down550 ) ,.TP42D1 ( pull_down582 )
     ,.TP34D1 ( pull_down614 ) ,.TP26D1 ( pull_down646 ) ,.TP18D1 ( pull_down678 )
     ,.TP50D0 ( pull_down551 ) ,.TP42D0 ( pull_down583 ) ,.TP34D0 ( pull_down615 )
     ,.TP26D0 ( pull_down647 ) ,.TP18D0 ( pull_down679 ) ,.TP41D3 ( pull_down584 )
     ,.TP33D3 ( pull_down616 ) ,.TP25D3 ( pull_down648 ) ,.TP17D3 ( pull_down680 )
     ,.TP41D2 ( pull_down585 ) ,.TP33D2 ( pull_down617 ) ,.TP25D2 ( pull_down649 )
     ,.TP17D2 ( pull_down681 ) ,.TP41D1 ( pull_down586 ) ,.TP33D1 ( pull_down618 )
     ,.TP25D1 ( pull_down650 ) ,.TP17D1 ( pull_down682 ) ,.TP41D0 ( pull_down587 )
     ,.TP33D0 ( pull_down619 ) ,.TP25D0 ( pull_down651 ) ,.TP17D0 ( pull_down683 )
     ,.TP40D3 ( pull_down588 ) ,.TP32D3 ( pull_down620 ) ,.TP24D3 ( pull_down652 )
     ,.TP16D3 ( pull_down684 ) ,.TP40D2 ( pull_down589 ) ,.TP32D2 ( pull_down621 )
     ,.TP24D2 ( pull_down653 ) ,.TP16D2 ( pull_down685 ) ,.TP40D1 ( pull_down590 )
     ,.TP32D1 ( pull_down622 ) ,.TP24D1 ( pull_down654 ) ,.TP16D1 ( pull_down686 )
     ,.TP40D0 ( pull_down591 ) ,.TP32D0 ( pull_down623 ) ,.TP24D0 ( pull_down655 )
     ,.TP16D0 ( pull_down687 ) ,.TP31D3 ( pull_down624 ) ,.TP23D3 ( pull_down656 )
     ,.TP15D3 ( pull_down688 ) ,.TP31D2 ( pull_down625 ) ,.TP23D2 ( pull_down657 )
     ,.TP15D2 ( pull_down689 ) ,.TP31D1 ( pull_down626 ) ,.TP23D1 ( pull_down658 )
     ,.TP15D1 ( pull_down690 ) ,.TP31D0 ( pull_down627 ) ,.TP23D0 ( pull_down659 )
     ,.TP15D0 ( pull_down691 ) ,.TP30D3 ( pull_down628 ) ,.TP22D3 ( pull_down660 )
     ,.TP14D3 ( pull_down692 ) ,.TP30D2 ( pull_down629 ) ,.TP22D2 ( pull_down661 )
     ,.TP14D2 ( pull_down693 ) ,.TP30D1 ( pull_down630 ) ,.TP22D1 ( pull_down662 )
     ,.TP14D1 ( pull_down694 ) ,.TP30D0 ( pull_down631 ) ,.TP22D0 ( pull_down663 )
     ,.TP14D0 ( pull_down695 ) ,.TP21D3 ( pull_down664 ) ,.TP13D3 ( pull_down696 )
     ,.TP21D2 ( pull_down665 ) ,.TP13D2 ( pull_down697 ) ,.TP21D1 ( pull_down666 )
     ,.TP13D1 ( pull_down698 ) ,.TP21D0 ( pull_down667 ) ,.TP13D0 ( pull_down699 )
     ,.TP20D3 ( pull_down668 ) ,.TP12D3 ( pull_down700 ) ,.TP20D2 ( pull_down669 )
     ,.TP12D2 ( pull_down701 ) ,.TP20D1 ( pull_down670 ) ,.TP12D1 ( pull_down702 )
     ,.TP20D0 ( pull_down671 ) ,.TP12D0 ( pull_down703 ) ,.TP11D3 ( pull_down704 )
     ,.TP11D2 ( pull_down705 ) ,.TP11D1 ( pull_down706 ) ,.TP11D0 ( pull_down707 )
     ,.TP10D3 ( pull_down708 ) ,.TP10D2 ( pull_down709 ) ,.TP10D1 ( pull_down710 )
     ,.TP10D0 ( pull_down711 ) ,.TP9D3 ( pull_down712 ) ,.TP9D2 ( pull_down713 )
     ,.TP9D1 ( pull_down714 ) ,.TP9D0 ( pull_down715 ) ,.TP8D3 ( pull_down716 )
     ,.TP8D2 ( pull_down717 ) ,.TP8D1 ( pull_down718 ) ,.TP8D0 ( pull_down719 )
     ,.TP7D3 ( pull_down720 ) ,.TP7D2 ( pull_down721 ) ,.TP7D1 ( pull_down722 )
     ,.TP7D0 ( pull_down723 ) ,.TP6D3 ( pull_down724 ) ,.TP6D2 ( pull_down725 )
     ,.TP6D1 ( pull_down726 ) ,.TP6D0 ( pull_down727 ) ,.TP5D3 ( pull_down728 )
     ,.TP5D2 ( pull_down729 ) ,.TP5D1 ( pull_down730 ) ,.TP5D0 ( pull_down731 )
     ,.TP4D3 ( pull_down732 ) ,.TP4D2 ( pull_down733 ) ,.TP4D1 ( pull_down734 )
     ,.TP4D0 ( pull_down735 ) ,.TP3D3 ( pull_down736 ) ,.TP3D2 ( pull_down737 )
     ,.TP3D1 ( pull_down738 ) ,.TP3D0 ( pull_down739 ) ,.TP2D3 ( pull_down740 )
     ,.TP2D2 ( pull_down741 ) ,.TP2D1 ( pull_down742 ) ,.TP2D0 ( pull_down743 )
     ,.TP1D3 ( pull_down744 ) ,.TP1D2 ( pull_down745 ) ,.TP1D1 ( pull_down746 )
     ,.TP1D0 ( pull_down747 ) ,.CLK30MHZ ( CLK30MHZ ) ,.EROMRDB ( EROMRDB )
     ,.EROMCSB ( EROMCSB ) ,.EROMPA2 ( EROMPA2 ) ,.EROMCLK ( EROMCLK )
     ,.EROMPA17 ( EROMPA17 ) ,.EROMPA16 ( EROMPA16 ) ,.EROMPA15 ( EROMPA15 )
     ,.EROMPA14 ( EROMPA14 ) ,.EROMPA13 ( EROMPA13 ) ,.EROMPA12 ( EROMPA12 )
     ,.EROMPA11 ( EROMPA11 ) ,.EROMPA10 ( EROMPA10 ) ,.EROMPA9 ( EROMPA9 )
     ,.EROMPD3 ( EROMPD3 ) ,.EROMPA8 ( EROMPA8 ) ,.EROMPD2 ( EROMPD2 )
     ,.EROMPA7 ( EROMPA7 ) ,.EROMPD1 ( EROMPD1 ) ,.EROMPA6 ( EROMPA6 )
     ,.EROMPD0 ( EROMPD0 ) ,.EROMPA5 ( EROMPA5 ) ,.EROMPA4 ( EROMPA4 )
     ,.EROMPA3 ( EROMPA3 ) ,.EROMPA1 ( EROMPA1 ) ,.EROMPA0 ( EROMPA0 )
     ,.RDCLKP1_OUT ( RDCLKP1_OUT ) ,.EXA_OUT ( EXA_OUT ) ,.WWR_OUT ( WWR_OUT )
     ,.CER_OUT ( CER_OUT ) ,.SER_OUT ( SER_OUT ) ,.EXER_OUT ( EXER_OUT )
     ,.MRG00_OUT ( MRG00_OUT ) ,.MRG01_OUT ( MRG01_OUT ) ,.MRG10_OUT ( MRG10_OUT )
     ,.MRG11_OUT ( MRG11_OUT ) ,.MRG12_OUT ( MRG12_OUT ) ,.DIS_OUT ( DIS_OUT )
     ,.READ_OUT ( READ_OUT ) ,.FCLK_OUT ( FCLK_OUT ) ,.PROGI_OUT ( PROGI_OUT )
     ,.BFA_OUT ( BFA_OUT ) ,.EROMPD31 ( EROMPD31 ) ,.EROMPD23 ( EROMPD23 )
     ,.EROMPD15 ( EROMPD15 ) ,.EROMPD30 ( EROMPD30 ) ,.EROMPD22 ( EROMPD22 )
     ,.EROMPD14 ( EROMPD14 ) ,.EROMPD29 ( EROMPD29 ) ,.EROMPD28 ( EROMPD28 )
     ,.EROMPD27 ( EROMPD27 ) ,.EROMPD19 ( EROMPD19 ) ,.EROMPD26 ( EROMPD26 )
     ,.EROMPD18 ( EROMPD18 ) ,.EROMPD25 ( EROMPD25 ) ,.EROMPD17 ( EROMPD17 )
     ,.EROMPD24 ( EROMPD24 ) ,.EROMPD16 ( EROMPD16 ) ,.EROMPD21 ( EROMPD21 )
     ,.EROMPD13 ( EROMPD13 ) ,.EROMPD20 ( EROMPD20 ) ,.EROMPD12 ( EROMPD12 )
     ,.EROMPD11 ( EROMPD11 ) ,.EROMPD10 ( EROMPD10 ) ,.EROMPD9 ( EROMPD9 )
     ,.EROMPD8 ( EROMPD8 ) ,.EROMPD7 ( EROMPD7 ) ,.EROMPD6 ( EROMPD6 )
     ,.EROMPD5 ( EROMPD5 ) ,.EROMPD4 ( EROMPD4 ) ,.BTFLG ( BTFLG ) ,.TMSPMD ( TMSPMD )
     ,.TMBTSEL ( TMBTSEL ) ,.ICETMSPMD ( ICETMSPMD ) ,.ICETMBTSEL ( ICETMBTSEL )
     ,.RESB ( RESB ) ,.USBCLK ( USBCLK ) ,.USBRD_B ( USBRD_B ) ,.USBWR0_B ( USBWR0_B )
     ,.USBA21 ( USBA21 ) ,.USBA20 ( USBA20 ) ,.USBA19 ( USBA19 ) ,.USBA4 ( USBA4 )
     ,.USBA3 ( USBA3 ) ,.USBA2 ( USBA2 ) ,.USBWAIT_B ( USBWAIT_B ) ,.USBD15 ( USBD15 )
     ,.USBD14 ( USBD14 ) ,.USBD13 ( USBD13 ) ,.USBD12 ( USBD12 ) ,.USBD11 ( USBD11 )
     ,.USBD10 ( USBD10 ) ,.USBD9 ( USBD9 ) ,.USBD8 ( USBD8 ) ,.USBD7 ( USBD7 )
     ,.USBD6 ( USBD6 ) ,.USBD5 ( USBD5 ) ,.USBD4 ( USBD4 ) ,.USBD3 ( USBD3 )
     ,.USBD2 ( USBD2 ) ,.USBD1 ( USBD1 ) ,.USBD0 ( USBD0 ) ,.ICESYSRES_B ( ICESYSRES_B )
     ,.ICECPURES_B ( ICECPURES_B ) ,.RESET_B ( RESET_B ) ,.EVAOSCMCLK ( EVAOSCMCLK )
     ,.EVAOSCRCLK1 ( pull_down4 ) ,.EVAOSCRCLK2 ( pull_down5 ) ,.EVAOSCRCLK3 ( pull_down6 )
     ,.TMEMA16 ( TMEMA16 ) ,.TMEMA15 ( TMEMA15 ) ,.TMEMA13 ( TMEMA13 )
     ,.TMEMA12 ( TMEMA12 ) ,.TMEMA11 ( TMEMA11 ) ,.TMEMA10 ( TMEMA10 )
     ,.TMEMA9 ( TMEMA9 ) ,.TMEMD3 ( TMEMD3 ) ,.TMEMA8 ( TMEMA8 ) ,.TMEMD2 ( TMEMD2 )
     ,.TMEMA7 ( TMEMA7 ) ,.TMEMD1 ( TMEMD1 ) ,.TMEMA6 ( TMEMA6 ) ,.TMEMD0 ( TMEMD0 )
     ,.TMEMA5 ( TMEMA5 ) ,.TMEMA4 ( TMEMA4 ) ,.TMEMA3 ( TMEMA3 ) ,.TMEMA2 ( TMEMA2 )
     ,.TMEMA1 ( TMEMA1 ) ,.TMEMA0 ( TMEMA0 ) ,.TMEMCS_B ( TMEMCS_B ) ,.TMEMRD_B ( TMEMRD_B )
     ,.TMEMWR_B ( TMEMWR_B ) ,.TMEMCLK2 ( TMEMCLK2 ) ,.TMEMCLK1 ( TMEMCLK1 )
     ,.TMEMCLK0 ( TMEMCLK0 ) ,.TMEMD107 ( TMEMD107 ) ,.TMEMD106 ( TMEMD106 )
     ,.TMEMD105 ( TMEMD105 ) ,.TMEMD104 ( TMEMD104 ) ,.TMEMD103 ( TMEMD103 )
     ,.TMEMD102 ( TMEMD102 ) ,.TMEMD101 ( TMEMD101 ) ,.TMEMD100 ( TMEMD100 )
     ,.TMEMD99 ( TMEMD99 ) ,.TMEMD98 ( TMEMD98 ) ,.TMEMD97 ( TMEMD97 )
     ,.TMEMD89 ( TMEMD89 ) ,.TMEMD96 ( TMEMD96 ) ,.TMEMD88 ( TMEMD88 )
     ,.TMEMD95 ( TMEMD95 ) ,.TMEMD87 ( TMEMD87 ) ,.TMEMD79 ( TMEMD79 )
     ,.TMEMD94 ( TMEMD94 ) ,.TMEMD86 ( TMEMD86 ) ,.TMEMD78 ( TMEMD78 )
     ,.TMEMD93 ( TMEMD93 ) ,.TMEMD85 ( TMEMD85 ) ,.TMEMD77 ( TMEMD77 )
     ,.TMEMD69 ( TMEMD69 ) ,.TMEMD92 ( TMEMD92 ) ,.TMEMD84 ( TMEMD84 )
     ,.TMEMD76 ( TMEMD76 ) ,.TMEMD68 ( TMEMD68 ) ,.TMEMD91 ( TMEMD91 )
     ,.TMEMD83 ( TMEMD83 ) ,.TMEMD75 ( TMEMD75 ) ,.TMEMD67 ( TMEMD67 )
     ,.TMEMD59 ( TMEMD59 ) ,.TMEMD90 ( TMEMD90 ) ,.TMEMD82 ( TMEMD82 )
     ,.TMEMD74 ( TMEMD74 ) ,.TMEMD66 ( TMEMD66 ) ,.TMEMD58 ( TMEMD58 )
     ,.TMEMD81 ( TMEMD81 ) ,.TMEMD73 ( TMEMD73 ) ,.TMEMD65 ( TMEMD65 )
     ,.TMEMD57 ( TMEMD57 ) ,.TMEMD49 ( TMEMD49 ) ,.TMEMD80 ( TMEMD80 )
     ,.TMEMD72 ( TMEMD72 ) ,.TMEMD64 ( TMEMD64 ) ,.TMEMD56 ( TMEMD56 )
     ,.TMEMD48 ( TMEMD48 ) ,.TMEMD71 ( TMEMD71 ) ,.TMEMD63 ( TMEMD63 )
     ,.TMEMD55 ( TMEMD55 ) ,.TMEMD47 ( TMEMD47 ) ,.TMEMD39 ( TMEMD39 )
     ,.TMEMD70 ( TMEMD70 ) ,.TMEMD62 ( TMEMD62 ) ,.TMEMD54 ( TMEMD54 )
     ,.TMEMD46 ( TMEMD46 ) ,.TMEMD38 ( TMEMD38 ) ,.TMEMD61 ( TMEMD61 )
     ,.TMEMD53 ( TMEMD53 ) ,.TMEMD45 ( TMEMD45 ) ,.TMEMD37 ( TMEMD37 )
     ,.TMEMD29 ( TMEMD29 ) ,.TMEMD60 ( TMEMD60 ) ,.TMEMD52 ( TMEMD52 )
     ,.TMEMD44 ( TMEMD44 ) ,.TMEMD36 ( TMEMD36 ) ,.TMEMD28 ( TMEMD28 )
     ,.TMEMD51 ( TMEMD51 ) ,.TMEMD43 ( TMEMD43 ) ,.TMEMD35 ( TMEMD35 )
     ,.TMEMD27 ( TMEMD27 ) ,.TMEMD19 ( TMEMD19 ) ,.TMEMD50 ( TMEMD50 )
     ,.TMEMD42 ( TMEMD42 ) ,.TMEMD34 ( TMEMD34 ) ,.TMEMD26 ( TMEMD26 )
     ,.TMEMD18 ( TMEMD18 ) ,.TMEMD41 ( TMEMD41 ) ,.TMEMD33 ( TMEMD33 )
     ,.TMEMD25 ( TMEMD25 ) ,.TMEMD17 ( TMEMD17 ) ,.TMEMD40 ( TMEMD40 )
     ,.TMEMD32 ( TMEMD32 ) ,.TMEMD24 ( TMEMD24 ) ,.TMEMD16 ( TMEMD16 )
     ,.TMEMD31 ( TMEMD31 ) ,.TMEMD23 ( TMEMD23 ) ,.TMEMD15 ( TMEMD15 )
     ,.TMEMD30 ( TMEMD30 ) ,.TMEMD22 ( TMEMD22 ) ,.TMEMD14 ( TMEMD14 )
     ,.TMEMD21 ( TMEMD21 ) ,.TMEMD13 ( TMEMD13 ) ,.TMEMD20 ( TMEMD20 )
     ,.TMEMD12 ( TMEMD12 ) ,.TMEMD11 ( TMEMD11 ) ,.TMEMD10 ( TMEMD10 )
     ,.TMEMD9 ( TMEMD9 ) ,.TMEMD8 ( TMEMD8 ) ,.TMEMD7 ( TMEMD7 ) ,.TMEMD6 ( TMEMD6 )
     ,.TMEMD5 ( TMEMD5 ) ,.TMEMD4 ( TMEMD4 ) ,.TCCONNECT_B ( TCCONNECT_B )
     ,.EACONNECT_B ( EACONNECT_B ) ,.TVDDON ( TVDDON ) ,.TVDDSEL ( TVDDSEL )
     ,.LEDTVDD_B ( LEDTVDD_B ) ,.LEDCLOCK_B ( LEDCLOCK_B ) ,.LEDRUN_B ( LEDRUN_B )
     ,.LEDRESET_B ( LEDRESET_B ) ,.LEDSTANDBY_B ( LEDSTANDBY_B ) ,.LEDWAIT_B ( LEDWAIT_B )
     ,.DCE0 ( DCE0 ) ,.DCLKSEL1 ( DCLKSEL1 ) ,.DCER ( DCER ) ,.DSER ( DSER )
     ,.DWWR ( DWWR ) ,.DWED ( DWED ) ,.DMRG00 ( DMRG00 ) ,.DMRG01 ( DMRG01 )
     ,.DMRG10 ( DMRG10 ) ,.DMRG11 ( DMRG11 ) ,.DMRG12 ( DMRG12 ) ,.DREAD ( DREAD )
     ,.AF19 ( AF19 ) ,.AF18 ( AF18 ) ,.AF17 ( AF17 ) ,.DA13 ( DA13 ) ,.AF16 ( AF16 )
     ,.DA12 ( DA12 ) ,.AF15 ( AF15 ) ,.DA11 ( DA11 ) ,.AF14 ( AF14 ) ,.DA10 ( DA10 )
     ,.AF13 ( AF13 ) ,.AF12 ( AF12 ) ,.AF11 ( AF11 ) ,.AF10 ( AF10 ) ,.AF9 ( AF9 )
     ,.DA7 ( DA7 ) ,.AF8 ( AF8 ) ,.DA6 ( DA6 ) ,.AF5 ( AF5 ) ,.DA3 ( DA3 )
     ,.AF4 ( AF4 ) ,.DA2 ( DA2 ) ,.AF3 ( AF3 ) ,.DA1 ( DA1 ) ,.AF2 ( AF2 )
     ,.DA0 ( DA0 ) ,.AF1 ( AF1 ) ,.AF0 ( AF0 ) ,.DRDCLK ( DRDCLK ) ,.DRDCLKC1 ( DRDCLKC1 )
     ,.DA9 ( DA9 ) ,.DA8 ( DA8 ) ,.DRO11 ( DRO011 ) ,.DRO10 ( DRO010 )
     ,.DRO9 ( DRO09 ) ,.DRO8 ( DRO08 ) ,.DRO7 ( DRO07 ) ,.DRO6 ( DRO06 )
     ,.DRO5 ( DRO05 ) ,.DRO4 ( DRO04 ) ,.DRO3 ( DRO03 ) ,.DRO2 ( DRO02 )
     ,.DRO1 ( DRO01 ) ,.DRO0 ( DRO00 ) ,.DDIS_OUT ( DDIS_OUT ) ,.DRDCLKP1_OUT ( DRDCLKP1_OUT )
     ,.DWWR_OUT ( DWWR_OUT ) ,.DCER_OUT ( DCER_OUT ) ,.DSER_OUT ( DSER_OUT )
     ,.DMRG00_OUT ( DMRG00_OUT ) ,.DMRG01_OUT ( DMRG01_OUT ) ,.DMRG10_OUT ( DMRG10_OUT )
     ,.DMRG11_OUT ( DMRG11_OUT ) ,.DMRG12_OUT ( DMRG12_OUT ) ,.DREAD_OUT ( DREAD_OUT )
     ,.DFCLK_OUT ( DFCLK_OUT ) ,.SLDFLASH ( SLDFLASH )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/_ice/_macro/_eva/_kx4/_056/port_iobuf.v
  port_iobuf port_iobuf (
    .P00ENI ( P00ENI ) ,.P00DIN ( P00DIN ) ,.P00ENO ( P00ENO ) ,.P00DOUT ( P00DOUT )
     ,.P00 ( P00 ) ,.P00PUON ( P00PUON ) ,.P00PUONOUT ( P00PUONOUT ) ,.P01ENI ( P01ENI )
     ,.P01DIN ( P01DIN ) ,.P01ENO ( P01ENO ) ,.P01DOUT ( P01DOUT ) ,.P01 ( P01 )
     ,.P01SELIN ( P01SELIN ) ,.PTTL01 ( P01 ) ,.P01PUON ( P01PUON ) ,.P01PUONOUT ( P01PUONOUT )
     ,.P02ENI ( P02ENI ) ,.P10ENI ( P10ENI ) ,.P02DIN ( P02DIN ) ,.P10DIN ( P10DIN )
     ,.P02ENO ( P02ENO ) ,.P10ENO ( P10ENO ) ,.P02DOUT ( P02DOUT ) ,.P10DOUT ( P10DOUT )
     ,.P02 ( P02 ) ,.P10 ( P10 ) ,.P02PUON ( P02PUON ) ,.P10PUON ( P10PUON )
     ,.P02PUONOUT ( P02PUONOUT ) ,.P10PUONOUT ( P10PUONOUT ) ,.P03ENI ( P03ENI )
     ,.P11ENI ( P11ENI ) ,.P03DIN ( P03DIN ) ,.P11DIN ( P11DIN ) ,.P03ENO ( P03ENO )
     ,.P11ENO ( P11ENO ) ,.P03DOUT ( P03DOUT ) ,.P11DOUT ( P11DOUT ) ,.P03 ( P03 )
     ,.P11 ( P11 ) ,.P03SELIN ( P03SELIN ) ,.P11SELIN ( P11SELIN ) ,.PTTL03 ( PTTL03 )
     ,.PTTL11 ( PTTL11 ) ,.P03PUON ( P03PUON ) ,.P11PUON ( P11PUON ) ,.P03PUONOUT ( P03PUONOUT )
     ,.P11PUONOUT ( P11PUONOUT ) ,.P04ENI ( P04ENI ) ,.P12ENI ( P12ENI )
     ,.P20ENI ( P20ENI ) ,.P04DIN ( P04DIN ) ,.P12DIN ( P12DIN ) ,.P20DIN ( P20DIN )
     ,.P04ENO ( P04ENO ) ,.P12ENO ( P12ENO ) ,.P20ENO ( P20ENO ) ,.P04DOUT ( P04DOUT )
     ,.P12DOUT ( P12DOUT ) ,.P20DOUT ( P20DOUT ) ,.P04 ( P04 ) ,.P12 ( P12 )
     ,.P20 ( P20 ) ,.P04SELIN ( P04SELIN ) ,.PTTL04 ( PTTL04 ) ,.P04PUON ( P04PUON )
     ,.P12PUON ( P12PUON ) ,.P04PUONOUT ( P04PUONOUT ) ,.P12PUONOUT ( P12PUONOUT )
     ,.P05ENI ( P05ENI ) ,.P13ENI ( P13ENI ) ,.P21ENI ( P21ENI ) ,.P05DIN ( P05DIN )
     ,.P13DIN ( P13DIN ) ,.P21DIN ( P21DIN ) ,.P05ENO ( P05ENO ) ,.P13ENO ( P13ENO )
     ,.P21ENO ( P21ENO ) ,.P05DOUT ( P05DOUT ) ,.P13DOUT ( P13DOUT ) ,.P21DOUT ( P21DOUT )
     ,.P05 ( P05 ) ,.P13 ( P13 ) ,.P21 ( P21 ) ,.AP1 ( AP1 ) ,.P05PUON ( P05PUON )
     ,.P13PUON ( P13PUON ) ,.P05PUONOUT ( P05PUONOUT ) ,.P13PUONOUT ( P13PUONOUT )
     ,.P06ENI ( P06ENI ) ,.P14ENI ( P14ENI ) ,.P22ENI ( P22ENI ) ,.P30ENI ( P30ENI )
     ,.P06DIN ( P06DIN ) ,.P14DIN ( P14DIN ) ,.P22DIN ( P22DIN ) ,.P30DIN ( P30DIN )
     ,.P06ENO ( P06ENO ) ,.P14ENO ( P14ENO ) ,.P22ENO ( P22ENO ) ,.P30ENO ( P30ENO )
     ,.P06DOUT ( P06DOUT ) ,.P14DOUT ( P14DOUT ) ,.P22DOUT ( P22DOUT )
     ,.P30DOUT ( P30DOUT ) ,.P06 ( P06 ) ,.P14 ( P14 ) ,.P22 ( P22 ) ,.P30 ( P30 )
     ,.AP2 ( AP2 ) ,.P06PUON ( P06PUON ) ,.P14PUON ( P14PUON ) ,.P30PUON ( P30PUON )
     ,.P06PUONOUT ( P06PUONOUT ) ,.P14PUONOUT ( P14PUONOUT ) ,.P30PUONOUT ( P30PUONOUT )
     ,.P10SELIN ( P10SELIN ) ,.PTTL10 ( PTTL10 ) ,.P13SELIN ( P13SELIN )
     ,.PTTL13 ( PTTL13 ) ,.P14SELIN ( P14SELIN ) ,.PTTL14 ( PTTL14 ) ,.P15ENI ( P15ENI )
     ,.P23ENI ( P23ENI ) ,.P31ENI ( P31ENI ) ,.P15DIN ( P15DIN ) ,.P23DIN ( P23DIN )
     ,.P31DIN ( P31DIN ) ,.P15ENO ( P15ENO ) ,.P23ENO ( P23ENO ) ,.P31ENO ( P31ENO )
     ,.P15DOUT ( P15DOUT ) ,.P23DOUT ( P23DOUT ) ,.P31DOUT ( P31DOUT )
     ,.P15 ( P15 ) ,.P23 ( P23 ) ,.P31 ( P31 ) ,.AP3 ( AP3 ) ,.P15SELIN ( P15SELIN )
     ,.PTTL15 ( PTTL15 ) ,.P15PUON ( P15PUON ) ,.P31PUON ( P31PUON ) ,.P15PUONOUT ( P15PUONOUT )
     ,.P31PUONOUT ( P31PUONOUT ) ,.P16ENI ( P16ENI ) ,.P24ENI ( P24ENI )
     ,.P40ENI ( P40ENI ) ,.P16DIN ( P16DIN ) ,.P24DIN ( P24DIN ) ,.P40DIN ( P40DIN )
     ,.P16ENO ( P16ENO ) ,.P24ENO ( P24ENO ) ,.P40ENO ( P40ENO ) ,.P16DOUT ( P16DOUT )
     ,.P24DOUT ( P24DOUT ) ,.P40DOUT ( P40DOUT ) ,.P16 ( P16 ) ,.P24 ( P24 )
     ,.P40 ( P40 ) ,.AP4 ( AP4 ) ,.P16SELIN ( P16SELIN ) ,.PTTL16 ( PTTL16 )
     ,.P16PUON ( P16PUON ) ,.P40PUON ( P40PUON ) ,.P16PUONOUT ( P16PUONOUT )
     ,.P40PUONOUT ( P40PUONOUT ) ,.P17ENI ( P17ENI ) ,.P25ENI ( P25ENI )
     ,.P41ENI ( P41ENI ) ,.P17DIN ( P17DIN ) ,.P25DIN ( P25DIN ) ,.P41DIN ( P41DIN )
     ,.P17ENO ( P17ENO ) ,.P25ENO ( P25ENO ) ,.P41ENO ( P41ENO ) ,.P17DOUT ( P17DOUT )
     ,.P25DOUT ( P25DOUT ) ,.P41DOUT ( P41DOUT ) ,.P17 ( P17 ) ,.P25 ( P25 )
     ,.P41 ( P41 ) ,.AP5 ( AP5 ) ,.P17SELIN ( P17SELIN ) ,.PTTL17 ( PTTL17 )
     ,.P17PUON ( P17PUON ) ,.P41PUON ( P41PUON ) ,.P17PUONOUT ( P17PUONOUT )
     ,.P41PUONOUT ( P41PUONOUT ) ,.P26ENI ( P26ENI ) ,.P42ENI ( P42ENI )
     ,.P50ENI ( P50ENI ) ,.P26DIN ( P26DIN ) ,.P42DIN ( P42DIN ) ,.P50DIN ( P50DIN )
     ,.P26ENO ( P26ENO ) ,.P42ENO ( P42ENO ) ,.P50ENO ( P50ENO ) ,.P26DOUT ( P26DOUT )
     ,.P42DOUT ( P42DOUT ) ,.P50DOUT ( P50DOUT ) ,.P26 ( P26 ) ,.P42 ( P42 )
     ,.P50 ( P50 ) ,.AP6 ( AP6 ) ,.P27ENI ( P27ENI ) ,.P43ENI ( P43ENI )
     ,.P51ENI ( P51ENI ) ,.P27DIN ( P27DIN ) ,.P43DIN ( P43DIN ) ,.P51DIN ( P51DIN )
     ,.P27ENO ( P27ENO ) ,.P43ENO ( P43ENO ) ,.P51ENO ( P51ENO ) ,.P27DOUT ( P27DOUT )
     ,.P43DOUT ( P43DOUT ) ,.P51DOUT ( P51DOUT ) ,.P27 ( P27 ) ,.P43 ( P43 )
     ,.P51 ( P51 ) ,.AP7 ( AP7 ) ,.P42PUON ( P42PUON ) ,.P50PUON ( P50PUON )
     ,.P42PUONOUT ( P42PUONOUT ) ,.P50PUONOUT ( P50PUONOUT ) ,.P43PUON ( P43PUON )
     ,.P51PUON ( P51PUON ) ,.P43PUONOUT ( P43PUONOUT ) ,.P51PUONOUT ( P51PUONOUT )
     ,.P52ENI ( P52ENI ) ,.P60ENI ( P60ENI ) ,.P52DIN ( P52DIN ) ,.P60DIN ( P60DIN )
     ,.P52ENO ( P52ENO ) ,.P60ENO ( P60ENO ) ,.P52DOUT ( P52DOUT ) ,.P60DOUT ( P60DOUT )
     ,.P52 ( P52 ) ,.P60 ( P60 ) ,.AP8 ( AP8 ) ,.P52PUON ( P52PUON ) ,.P52PUONOUT ( P52PUONOUT )
     ,.P53ENI ( P53ENI ) ,.P61ENI ( P61ENI ) ,.DGEN01 ( DGEN01 ) ,.P53DIN ( P53DIN )
     ,.P61DIN ( P61DIN ) ,.P53ENO ( P53ENO ) ,.P61ENO ( P61ENO ) ,.DGEN07 ( DGEN07 )
     ,.P53DOUT ( P53DOUT ) ,.P61DOUT ( P61DOUT ) ,.P53 ( P53 ) ,.P61 ( P61 )
     ,.AP9 ( AP9 ) ,.P53PUON ( P53PUON ) ,.P53PUONOUT ( P53PUONOUT ) ,.P54ENI ( P54ENI )
     ,.P62ENI ( P62ENI ) ,.P70ENI ( P70ENI ) ,.P54DIN ( P54DIN ) ,.P62DIN ( P62DIN )
     ,.P70DIN ( P70DIN ) ,.DGEN00 ( DGEN00 ) ,.P54ENO ( P54ENO ) ,.P62ENO ( P62ENO )
     ,.P70ENO ( P70ENO ) ,.P54DOUT ( P54DOUT ) ,.P62DOUT ( P62DOUT ) ,.P70DOUT ( P70DOUT )
     ,.P54 ( P54 ) ,.P62 ( P62 ) ,.P70 ( P70 ) ,.P54PUON ( P54PUON ) ,.P70PUON ( P70PUON )
     ,.P54PUONOUT ( P54PUONOUT ) ,.P70PUONOUT ( P70PUONOUT ) ,.P55ENI ( P55ENI )
     ,.P63ENI ( P63ENI ) ,.P71ENI ( P71ENI ) ,.P55DIN ( P55DIN ) ,.P63DIN ( P63DIN )
     ,.P71DIN ( P71DIN ) ,.P55ENO ( P55ENO ) ,.P63ENO ( P63ENO ) ,.P71ENO ( P71ENO )
     ,.P55DOUT ( P55DOUT ) ,.P63DOUT ( P63DOUT ) ,.P71DOUT ( P71DOUT )
     ,.P55SELIN ( P55SELIN ) ,.P55 ( P55 ) ,.P63 ( P63 ) ,.P71 ( P71 )
     ,.PTTL55 ( P55 ) ,.P55PUON ( P55PUON ) ,.P71PUON ( P71PUON ) ,.P55PUONOUT ( P55PUONOUT )
     ,.P71PUONOUT ( P71PUONOUT ) ,.P72ENI ( P72ENI ) ,.P72DIN ( P72DIN )
     ,.P72ENO ( P72ENO ) ,.P72DOUT ( P72DOUT ) ,.P72 ( P72 ) ,.P72PUON ( P72PUON )
     ,.P72PUONOUT ( P72PUONOUT ) ,.P73ENI ( P73ENI ) ,.P73DIN ( P73DIN )
     ,.P73ENO ( P73ENO ) ,.P73DOUT ( P73DOUT ) ,.P73 ( P73 ) ,.P73PUON ( P73PUON )
     ,.P73PUONOUT ( P73PUONOUT ) ,.P74ENI ( P74ENI ) ,.P74DIN ( P74DIN )
     ,.P74ENO ( P74ENO ) ,.P74DOUT ( P74DOUT ) ,.P74 ( P74 ) ,.P74PUON ( P74PUON )
     ,.P74PUONOUT ( P74PUONOUT ) ,.P75ENI ( P75ENI ) ,.P75DIN ( P75DIN )
     ,.P75ENO ( P75ENO ) ,.P75DOUT ( P75DOUT ) ,.P75 ( P75 ) ,.P75PUON ( P75PUON )
     ,.P75PUONOUT ( P75PUONOUT ) ,.P76ENI ( P76ENI ) ,.P76DIN ( P76DIN )
     ,.P76ENO ( P76ENO ) ,.P76DOUT ( P76DOUT ) ,.P76 ( P76 ) ,.P76PUON ( P76PUON )
     ,.P76PUONOUT ( P76PUONOUT ) ,.P77ENI ( P77ENI ) ,.P77DIN ( P77DIN )
     ,.P77ENO ( P77ENO ) ,.P77DOUT ( P77DOUT ) ,.P77 ( P77 ) ,.P77PUON ( P77PUON )
     ,.P77PUONOUT ( P77PUONOUT ) ,.P120ENI ( P120ENI ) ,.P120DIN ( P120DIN )
     ,.P120ENO ( P120ENO ) ,.P120DOUT ( P120DOUT ) ,.P120 ( P120 ) ,.P120PUON ( P120PUON )
     ,.P120PUONOUT ( P120PUONOUT ) ,.P130ENO ( P130ENO ) ,.P130DOUT ( P130DOUT )
     ,.P130 ( P130 ) ,.AP10 ( AP10 ) ,.P137ENI ( P137ENI ) ,.P137DIN ( P137DIN )
     ,.P137 ( P137 ) ,.AP17 ( AP17 ) ,.AP25 ( AP25 ) ,.AP33 ( AP33 ) ,.AP41 ( AP41 )
     ,.P140ENI ( P140ENI ) ,.P140DIN ( P140DIN ) ,.P140ENO ( P140ENO )
     ,.P140DOUT ( P140DOUT ) ,.P140 ( P140 ) ,.AP12 ( AP12 ) ,.AP20 ( AP20 )
     ,.P140PUON ( P140PUON ) ,.P140PUONOUT ( P140PUONOUT ) ,.P141ENI ( P141ENI )
     ,.P141DIN ( P141DIN ) ,.P141ENO ( P141ENO ) ,.P141DOUT ( P141DOUT )
     ,.P141 ( P141 ) ,.AP13 ( AP13 ) ,.AP21 ( AP21 ) ,.P141PUON ( P141PUON )
     ,.P141PUONOUT ( P141PUONOUT ) ,.P146ENI ( P146ENI ) ,.P146DIN ( P146DIN )
     ,.P146ENO ( P146ENO ) ,.P146DOUT ( P146DOUT ) ,.P146 ( P146 ) ,.AP18 ( AP18 )
     ,.AP26 ( AP26 ) ,.AP34 ( AP34 ) ,.AP42 ( AP42 ) ,.AP50 ( AP50 ) ,.P146PUON ( P146PUON )
     ,.P146PUONOUT ( P146PUONOUT ) ,.P147ENI ( P147ENI ) ,.P147DIN ( P147DIN )
     ,.P147ENO ( P147ENO ) ,.P147DOUT ( P147DOUT ) ,.P147 ( P147 ) ,.AP19 ( AP19 )
     ,.AP27 ( AP27 ) ,.AP35 ( AP35 ) ,.AP43 ( AP43 ) ,.AP51 ( AP51 ) ,.P147PUON ( P147PUON )
     ,.P147PUONOUT ( P147PUONOUT ) ,.DGEN02 ( DGEN02 ) ,.DGEN03 ( DGEN03 )
     ,.DGEN04 ( DGEN04 ) ,.DGEN05 ( DGEN05 ) ,.DGEN06 ( DGEN06 ) ,.PORTEN_B0 ( PORTEN_B0 )
     ,.PORTEN_B1 ( PORTEN_B1 ) ,.PORTEN_B2 ( PORTEN_B2 ) ,.PORTEN_B3 ( PORTEN_B3 )
     ,.PORTEN_B4 ( PORTEN_B4 ) ,.PORTEN_B5 ( PORTEN_B5 ) ,.PORTEN_B6 ( PORTEN_B6 )
     ,.PORTEN_B7 ( PORTEN_B7 ) ,.PORTEN_B8 ( PORTEN_B8 ) ,.PORTEN_B9 ( PORTEN_B9 )
     ,.PORTEN_B10 ( PORTEN_B10 ) ,.PORTEN_B11 ( PORTEN_B11 ) ,.ADVSELMOD0_I ( ADVSELMOD0_I )
     ,.ADVSELMOD1_I ( ADVSELMOD1_I ) ,.EMVDDSEL_B ( EMVDDSEL_B ) ,.ADVSELMOD ( ADVSELMOD )
     ,.STOPZ ( STOPZ ) ,.RESFB5V ( RESFB5V ) ,.AP11 ( AP11 ) ,.AP14 ( AP14 )
     ,.AP22 ( AP22 ) ,.AP30 ( AP30 ) ,.AP15 ( AP15 ) ,.AP23 ( AP23 ) ,.AP31 ( AP31 )
     ,.AP16 ( AP16 ) ,.AP24 ( AP24 ) ,.AP32 ( AP32 ) ,.AP40 ( AP40 ) ,.AP28 ( AP28 )
     ,.AP36 ( AP36 ) ,.AP44 ( AP44 ) ,.AP52 ( AP52 ) ,.AP60 ( AP60 ) ,.AP29 ( AP29 )
     ,.AP37 ( AP37 ) ,.AP45 ( AP45 ) ,.AP53 ( AP53 ) ,.AP61 ( AP61 ) ,.AP38 ( AP38 )
     ,.AP46 ( AP46 ) ,.AP54 ( AP54 ) ,.AP62 ( AP62 ) ,.AP39 ( AP39 ) ,.AP47 ( AP47 )
     ,.AP55 ( AP55 ) ,.AP63 ( AP63 ) ,.AP48 ( AP48 ) ,.AP56 ( AP56 ) ,.AP64 ( AP64 )
     ,.AP49 ( AP49 ) ,.AP57 ( AP57 ) ,.AP65 ( AP65 ) ,.AP58 ( AP58 ) ,.AP59 ( AP59 )
     ,.APIO1 ( APIO1 ) ,.APIO2 ( APIO2 ) ,.APIO3 ( APIO3 ) ,.APIO4 ( APIO4 )
     ,.APIO5 ( APIO5 ) ,.APIO6 ( APIO6 ) ,.APIO7 ( APIO7 ) ,.APIO8 ( APIO8 )
     ,.APIO9 ( APIO9 ) ,.APIO10 ( APIO10 ) ,.APIO11 ( APIO11 ) ,.APIO12 ( APIO12 )
     ,.APIO20 ( APIO20 ) ,.APIO13 ( APIO13 ) ,.APIO21 ( APIO21 ) ,.APIO14 ( APIO14 )
     ,.APIO22 ( APIO22 ) ,.APIO30 ( APIO30 ) ,.APIO15 ( APIO15 ) ,.APIO23 ( APIO23 )
     ,.APIO31 ( APIO31 ) ,.APIO16 ( APIO16 ) ,.APIO24 ( APIO24 ) ,.APIO32 ( APIO32 )
     ,.APIO40 ( APIO40 ) ,.APIO17 ( APIO17 ) ,.APIO25 ( APIO25 ) ,.APIO33 ( APIO33 )
     ,.APIO41 ( APIO41 ) ,.APIO18 ( APIO18 ) ,.APIO26 ( APIO26 ) ,.APIO34 ( APIO34 )
     ,.APIO42 ( APIO42 ) ,.APIO50 ( APIO50 ) ,.APIO19 ( APIO19 ) ,.APIO27 ( APIO27 )
     ,.APIO35 ( APIO35 ) ,.APIO43 ( APIO43 ) ,.APIO51 ( APIO51 ) ,.APIO28 ( APIO28 )
     ,.APIO36 ( APIO36 ) ,.APIO44 ( APIO44 ) ,.APIO52 ( APIO52 ) ,.APIO60 ( APIO60 )
     ,.APIO29 ( APIO29 ) ,.APIO37 ( APIO37 ) ,.APIO45 ( APIO45 ) ,.APIO53 ( APIO53 )
     ,.APIO61 ( APIO61 ) ,.APIO38 ( APIO38 ) ,.APIO46 ( APIO46 ) ,.APIO54 ( APIO54 )
     ,.APIO62 ( APIO62 ) ,.APIO39 ( APIO39 ) ,.APIO47 ( APIO47 ) ,.APIO55 ( APIO55 )
     ,.APIO63 ( APIO63 ) ,.APIO48 ( APIO48 ) ,.APIO56 ( APIO56 ) ,.APIO64 ( APIO64 )
     ,.APIO49 ( APIO49 ) ,.APIO57 ( APIO57 ) ,.APIO65 ( APIO65 ) ,.APIO58 ( APIO58 )
     ,.APIO59 ( APIO59 ) ,.PIO_ANALOG0 ( PIO_ANALOG0 ) ,.PIO_ANALOG1 ( PIO_ANALOG1 )
     ,.PIO_ANALOG2 ( PIO_ANALOG2 ) ,.PIO_ANALOG3 ( PIO_ANALOG3 ) ,.PIO_ANALOG4 ( PIO_ANALOG4 )
     ,.PIO_ANALOG5 ( PIO_ANALOG5 ) ,.PORTEN_B12 ( PORTEN_B12 ) ,.PORTEN_B20 ( PORTEN_B20 )
     ,.PORTEN_B13 ( PORTEN_B13 ) ,.PORTEN_B21 ( PORTEN_B21 ) ,.PORTEN_B14 ( PORTEN_B14 )
     ,.PORTEN_B22 ( PORTEN_B22 ) ,.PORTEN_B15 ( PORTEN_B15 ) ,.PORTEN_B23 ( PORTEN_B23 )
     ,.PORTEN_B16 ( PORTEN_B16 ) ,.PORTEN_B24 ( PORTEN_B24 ) ,.PORTEN_B17 ( PORTEN_B17 )
     ,.PORTEN_B25 ( PORTEN_B25 ) ,.PORTEN_B18 ( PORTEN_B18 ) ,.PORTEN_B26 ( PORTEN_B26 )
     ,.PORTEN_B19 ( PORTEN_B19 )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/_ice/_macro/_eva/_kx4/_056/puctl6.v
  PUCTL puctl (
    .CLK60MHZ ( CLK60MHZ ) ,.CPURSOUTB ( SYSRSOUTB ) ,.DIN000 ( pull_down33 )
     ,.DIN001 ( pull_down34 ) ,.DIN002 ( pull_down35 ) ,.DIN010 ( pull_down43 )
     ,.DIN003 ( pull_down36 ) ,.DIN011 ( pull_down44 ) ,.DIN004 ( pull_down37 )
     ,.DIN012 ( P30PUONOUT ) ,.DIN020 ( P76PUONOUT ) ,.DIN100 ( pull_down53 )
     ,.DIN005 ( pull_down38 ) ,.DIN013 ( P31PUONOUT ) ,.DIN021 ( P77PUONOUT )
     ,.DIN101 ( pull_down54 ) ,.DIN006 ( pull_down39 ) ,.DIN014 ( P70PUONOUT )
     ,.DIN030 ( pull_down51 ) ,.DIN102 ( pull_down55 ) ,.DIN110 ( pull_down63 )
     ,.DIN007 ( pull_down40 ) ,.DIN015 ( P71PUONOUT ) ,.DIN031 ( pull_down52 )
     ,.DIN103 ( pull_down56 ) ,.DIN111 ( pull_down64 ) ,.DIN008 ( pull_down41 )
     ,.DIN016 ( P72PUONOUT ) ,.DIN024 ( pull_down45 ) ,.DIN104 ( pull_down57 )
     ,.DIN112 ( pull_down65 ) ,.DIN120 ( pull_down73 ) ,.DIN200 ( pull_down83 )
     ,.DIN009 ( pull_down42 ) ,.DIN017 ( P73PUONOUT ) ,.DIN025 ( pull_down46 )
     ,.DIN105 ( pull_down58 ) ,.DIN113 ( pull_down66 ) ,.DIN121 ( pull_down74 )
     ,.DIN201 ( pull_down84 ) ,.DIN018 ( P74PUONOUT ) ,.DIN026 ( pull_down47 )
     ,.DIN106 ( pull_down59 ) ,.DIN114 ( pull_down67 ) ,.DIN130 ( pull_down81 )
     ,.DIN202 ( pull_down85 ) ,.DIN210 ( pull_down93 ) ,.DIN019 ( P75PUONOUT )
     ,.DIN027 ( pull_down48 ) ,.DIN107 ( pull_down60 ) ,.DIN115 ( pull_down68 )
     ,.DIN131 ( pull_down82 ) ,.DIN203 ( pull_down86 ) ,.DIN211 ( pull_down94 )
     ,.DIN028 ( pull_down49 ) ,.DIN108 ( pull_down61 ) ,.DIN116 ( pull_down69 )
     ,.DIN124 ( pull_down75 ) ,.DIN204 ( pull_down87 ) ,.DIN212 ( P10PUONOUT )
     ,.DIN220 ( pull_down95 ) ,.DIN300 ( pull_down105 ) ,.DIN029 ( pull_down50 )
     ,.DIN109 ( pull_down62 ) ,.DIN117 ( pull_down70 ) ,.DIN125 ( pull_down76 )
     ,.DIN205 ( pull_down88 ) ,.DIN213 ( P11PUONOUT ) ,.DIN221 ( pull_down96 )
     ,.DIN301 ( pull_down106 ) ,.DIN118 ( pull_down71 ) ,.DIN126 ( pull_down77 )
     ,.DIN206 ( pull_down89 ) ,.DIN214 ( P12PUONOUT ) ,.DIN230 ( pull_down103 )
     ,.DIN302 ( pull_down107 ) ,.DIN310 ( pull_down115 ) ,.DIN119 ( pull_down72 )
     ,.DIN127 ( pull_down78 ) ,.DIN207 ( pull_down90 ) ,.DIN215 ( P13PUONOUT )
     ,.DIN231 ( pull_down104 ) ,.DIN303 ( pull_down108 ) ,.DIN311 ( pull_down116 )
     ,.DIN128 ( pull_down79 ) ,.DIN208 ( pull_down91 ) ,.DIN216 ( P14PUONOUT )
     ,.DIN224 ( pull_down97 ) ,.DIN304 ( pull_down109 ) ,.DIN312 ( pull_down117 )
     ,.DIN320 ( pull_down121 ) ,.DIN400 ( pull_down125 ) ,.DIN129 ( pull_down80 )
     ,.DIN209 ( pull_down92 ) ,.DIN217 ( P15PUONOUT ) ,.DIN225 ( pull_down98 )
     ,.DIN305 ( pull_down110 ) ,.DIN313 ( P40PUONOUT ) ,.DIN321 ( pull_down122 )
     ,.DIN401 ( pull_down126 ) ,.DIN218 ( P16PUONOUT ) ,.DIN226 ( pull_down99 )
     ,.DIN306 ( pull_down111 ) ,.DIN314 ( P41PUONOUT ) ,.DIN330 ( pull_down123 )
     ,.DIN402 ( pull_down127 ) ,.DIN410 ( pull_down135 ) ,.DIN219 ( P17PUONOUT )
     ,.DIN227 ( pull_down100 ) ,.DIN307 ( pull_down112 ) ,.DIN315 ( P42PUONOUT )
     ,.DIN331 ( pull_down124 ) ,.DIN403 ( pull_down128 ) ,.DIN411 ( pull_down136 )
     ,.DIN228 ( pull_down101 ) ,.DIN308 ( pull_down113 ) ,.DIN316 ( P43PUONOUT )
     ,.DIN324 ( P50PUONOUT ) ,.DIN404 ( pull_down129 ) ,.DIN412 ( P00PUONOUT )
     ,.DIN420 ( pull_down140 ) ,.DIN500 ( pull_down147 ) ,.DIN229 ( pull_down102 )
     ,.DIN309 ( pull_down114 ) ,.DIN317 ( pull_down118 ) ,.DIN325 ( P51PUONOUT )
     ,.DIN405 ( pull_down130 ) ,.DIN413 ( P01PUONOUT ) ,.DIN421 ( pull_down141 )
     ,.DIN501 ( pull_down148 ) ,.DIN318 ( pull_down119 ) ,.DIN326 ( P52PUONOUT )
     ,.DIN406 ( pull_down131 ) ,.DIN414 ( pull_down137 ) ,.DIN430 ( P146PUONOUT )
     ,.DIN502 ( pull_down149 ) ,.DIN510 ( pull_down157 ) ,.DIN319 ( pull_down120 )
     ,.DIN327 ( P53PUONOUT ) ,.DIN407 ( pull_down132 ) ,.DIN415 ( pull_down138 )
     ,.DIN431 ( pull_down146 ) ,.DIN503 ( pull_down150 ) ,.DIN511 ( pull_down158 )
     ,.DIN328 ( P54PUONOUT ) ,.DIN408 ( pull_down133 ) ,.DIN416 ( P04PUONOUT )
     ,.DIN424 ( pull_down142 ) ,.DIN504 ( pull_down151 ) ,.DIN512 ( pull_down159 )
     ,.DIN520 ( pull_down162 ) ,.DIN329 ( P55PUONOUT ) ,.DIN409 ( pull_down134 )
     ,.DIN417 ( P05PUONOUT ) ,.DIN425 ( pull_down143 ) ,.DIN505 ( pull_down152 )
     ,.DIN513 ( pull_down160 ) ,.DIN521 ( pull_down163 ) ,.DIN418 ( P06PUONOUT )
     ,.DIN426 ( pull_down144 ) ,.DIN506 ( pull_down153 ) ,.DIN514 ( P02PUONOUT )
     ,.DIN530 ( pull_down170 ) ,.DIN419 ( pull_down139 ) ,.DIN427 ( pull_down145 )
     ,.DIN507 ( pull_down154 ) ,.DIN515 ( P03PUONOUT ) ,.DIN531 ( pull_down171 )
     ,.DIN428 ( P140PUONOUT ) ,.DIN508 ( pull_down155 ) ,.DIN516 ( P120PUONOUT )
     ,.DIN524 ( pull_down164 ) ,.DIN429 ( P141PUONOUT ) ,.DIN509 ( pull_down156 )
     ,.DIN517 ( P120PUONOUT ) ,.DIN525 ( pull_down165 ) ,.DIN518 ( P147PUONOUT )
     ,.DIN526 ( pull_down166 ) ,.DIN519 ( pull_down161 ) ,.DIN527 ( pull_down167 )
     ,.DIN528 ( pull_down168 ) ,.DIN529 ( pull_down169 ) ,.PSSC0L ( pull_up2 )
     ,.PPUP16 ( PPUP16 ) ,.PPUP24 ( PPUP24 ) ,.PSSC1L ( pull_down30 ) ,.PPUP18 ( PPUP18 )
     ,.PPUP26 ( PPUP26 ) ,.PSSC2L ( pull_up3 ) ,.PPUP28 ( PPUP28 ) ,.PSSC3L ( pull_down31 )
     ,.PSSC4L ( pull_down32 ) ,.PSSC5L ( pull_up4 ) ,.PPUP0 ( PPUP0 ) ,.PPUP1 ( PPUP1 )
     ,.PPUP2 ( PPUP2 ) ,.PPUP3 ( PPUP3 ) ,.PPUP4 ( PPUP4 ) ,.PPUP5 ( PPUP5 )
     ,.PPUP6 ( PPUP6 ) ,.PPUP7 ( PPUP7 ) ,.PPUP8 ( PPUP8 ) ,.PPUP9 ( PPUP9 )
     ,.PPUP10 ( PPUP10 ) ,.PPUP11 ( PPUP11 ) ,.PPUP12 ( PPUP12 ) ,.PPUP20 ( PPUP20 )
     ,.PPUP13 ( PPUP13 ) ,.PPUP21 ( PPUP21 ) ,.PPUP14 ( PPUP14 ) ,.PPUP30 ( PPUP30 )
     ,.PPUP15 ( PPUP15 ) ,.PPUP31 ( PPUP31 ) ,.PPUP17 ( PPUP17 ) ,.PPUP25 ( PPUP25 )
     ,.PPUP19 ( PPUP19 ) ,.PPUP27 ( PPUP27 ) ,.PPUP29 ( PPUP29 ) ,.PSSC0 ( PSSC0 )
     ,.PSSC1 ( PSSC1 ) ,.PSSC2 ( PSSC2 ) ,.PSSC3 ( PSSC3 ) ,.PSSC4 ( PSSC4 )
     ,.PSSC5 ( PSSC5 ) ,.PUPLE0 ( PUPLE0 ) ,.PUPLE1 ( PUPLE1 ) ,.PUPLE2 ( PUPLE2 )
     ,.PUPLE3 ( PUPLE3 ) ,.PUPLE4 ( PUPLE4 ) ,.PUPLE5 ( PUPLE5 )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/_ice/_macro/_eva/_kx4/_056/evatop_other.v
  evatop_other evatop_other (
    .ADDRTD144 ( ADDRTD144 ) ,.ADDRTD136 ( ADDRTD136 ) ,.ADDRTD128 ( ADDRTD128 )
     ,.ADDRTD143 ( ADDRTD143 ) ,.ADDRTD135 ( ADDRTD135 ) ,.ADDRTD127 ( ADDRTD127 )
     ,.ADDRTD119 ( ADDRTD119 ) ,.ADDRTD142 ( ADDRTD142 ) ,.ADDRTD134 ( ADDRTD134 )
     ,.ADDRTD126 ( ADDRTD126 ) ,.ADDRTD118 ( ADDRTD118 ) ,.ADDRTD141 ( ADDRTD141 )
     ,.ADDRTD133 ( ADDRTD133 ) ,.ADDRTD125 ( ADDRTD125 ) ,.ADDRTD117 ( ADDRTD117 )
     ,.ADDRTD109 ( ADDRTD109 ) ,.ADDRTD140 ( ADDRTD140 ) ,.ADDRTD132 ( ADDRTD132 )
     ,.ADDRTD124 ( ADDRTD124 ) ,.ADDRTD116 ( ADDRTD116 ) ,.ADDRTD108 ( ADDRTD108 )
     ,.ADDRTD139 ( ADDRTD139 ) ,.ADDRTD138 ( ADDRTD138 ) ,.ADDRTD137 ( ADDRTD137 )
     ,.ADDRTD129 ( ADDRTD129 ) ,.ADDRTD131 ( ADDRTD131 ) ,.ADDRTD123 ( ADDRTD123 )
     ,.ADDRTD115 ( ADDRTD115 ) ,.ADDRTD107 ( ADDRTD107 ) ,.ADDRTD130 ( ADDRTD130 )
     ,.ADDRTD122 ( ADDRTD122 ) ,.ADDRTD114 ( ADDRTD114 ) ,.ADDRTD106 ( ADDRTD106 )
     ,.ADDRTD121 ( ADDRTD121 ) ,.ADDRTD113 ( ADDRTD113 ) ,.ADDRTD105 ( ADDRTD105 )
     ,.ADDRTD120 ( ADDRTD120 ) ,.ADDRTD112 ( ADDRTD112 ) ,.ADDRTD104 ( ADDRTD104 )
     ,.ADDRTD111 ( ADDRTD111 ) ,.ADDRTD103 ( ADDRTD103 ) ,.ADDRTD110 ( ADDRTD110 )
     ,.ADDRTD102 ( ADDRTD102 ) ,.ADDRTD101 ( ADDRTD101 ) ,.ADDRTD100 ( ADDRTD100 )
     ,.ADDRTD99 ( ADDRTD99 ) ,.ADDRTD98 ( ADDRTD98 ) ,.ADDRTD97 ( ADDRTD97 )
     ,.ADDRTD89 ( ADDRTD89 ) ,.ADDRTD96 ( ADDRTD96 ) ,.ADDRTD88 ( ADDRTD88 )
     ,.ADDRTD95 ( ADDRTD95 ) ,.ADDRTD87 ( ADDRTD87 ) ,.ADDRTD79 ( ADDRTD79 )
     ,.ADDRTD94 ( ADDRTD94 ) ,.ADDRTD86 ( ADDRTD86 ) ,.ADDRTD78 ( ADDRTD78 )
     ,.ADDRTD93 ( ADDRTD93 ) ,.ADDRTD85 ( ADDRTD85 ) ,.ADDRTD77 ( ADDRTD77 )
     ,.ADDRTD69 ( ADDRTD69 ) ,.ADDRTD92 ( ADDRTD92 ) ,.ADDRTD84 ( ADDRTD84 )
     ,.ADDRTD76 ( ADDRTD76 ) ,.ADDRTD68 ( ADDRTD68 ) ,.ADDRTD91 ( ADDRTD91 )
     ,.ADDRTD83 ( ADDRTD83 ) ,.ADDRTD75 ( ADDRTD75 ) ,.ADDRTD67 ( ADDRTD67 )
     ,.ADDRTD59 ( ADDRTD59 ) ,.ADDRTD90 ( ADDRTD90 ) ,.ADDRTD82 ( ADDRTD82 )
     ,.ADDRTD74 ( ADDRTD74 ) ,.ADDRTD66 ( ADDRTD66 ) ,.ADDRTD58 ( ADDRTD58 )
     ,.ADDRTD81 ( ADDRTD81 ) ,.ADDRTD73 ( ADDRTD73 ) ,.ADDRTD65 ( ADDRTD65 )
     ,.ADDRTD57 ( ADDRTD57 ) ,.ADDRTD49 ( ADDRTD49 ) ,.ADDRTD80 ( ADDRTD80 )
     ,.ADDRTD72 ( ADDRTD72 ) ,.ADDRTD64 ( ADDRTD64 ) ,.ADDRTD56 ( ADDRTD56 )
     ,.ADDRTD48 ( ADDRTD48 ) ,.ADDRTD71 ( ADDRTD71 ) ,.ADDRTD63 ( ADDRTD63 )
     ,.ADDRTD55 ( ADDRTD55 ) ,.ADDRTD47 ( ADDRTD47 ) ,.ADDRTD39 ( ADDRTD39 )
     ,.ADDRTD70 ( ADDRTD70 ) ,.ADDRTD62 ( ADDRTD62 ) ,.ADDRTD54 ( ADDRTD54 )
     ,.ADDRTD46 ( ADDRTD46 ) ,.ADDRTD38 ( ADDRTD38 ) ,.ADDRTD61 ( ADDRTD61 )
     ,.ADDRTD53 ( ADDRTD53 ) ,.ADDRTD45 ( ADDRTD45 ) ,.ADDRTD37 ( ADDRTD37 )
     ,.ADDRTD29 ( ADDRTD29 ) ,.ADDRTD60 ( ADDRTD60 ) ,.ADDRTD52 ( ADDRTD52 )
     ,.ADDRTD44 ( ADDRTD44 ) ,.ADDRTD36 ( ADDRTD36 ) ,.ADDRTD28 ( ADDRTD28 )
     ,.ADDRTD51 ( ADDRTD51 ) ,.ADDRTD43 ( ADDRTD43 ) ,.ADDRTD35 ( ADDRTD35 )
     ,.ADDRTD27 ( ADDRTD27 ) ,.ADDRTD19 ( ADDRTD19 ) ,.ADDRTD50 ( ADDRTD50 )
     ,.ADDRTD42 ( ADDRTD42 ) ,.ADDRTD34 ( ADDRTD34 ) ,.ADDRTD26 ( ADDRTD26 )
     ,.ADDRTD18 ( ADDRTD18 ) ,.ADDRTD41 ( ADDRTD41 ) ,.ADDRTD33 ( ADDRTD33 )
     ,.ADDRTD25 ( ADDRTD25 ) ,.ADDRTD17 ( ADDRTD17 ) ,.ADDRTD40 ( ADDRTD40 )
     ,.ADDRTD32 ( ADDRTD32 ) ,.ADDRTD24 ( ADDRTD24 ) ,.ADDRTD16 ( ADDRTD16 )
     ,.ADDRTD31 ( ADDRTD31 ) ,.ADDRTD23 ( ADDRTD23 ) ,.ADDRTD15 ( ADDRTD15 )
     ,.ADDRTD30 ( ADDRTD30 ) ,.ADDRTD22 ( ADDRTD22 ) ,.ADDRTD14 ( ADDRTD14 )
     ,.ADDRTD21 ( ADDRTD21 ) ,.ADDRTD13 ( ADDRTD13 ) ,.ADDRTD20 ( ADDRTD20 )
     ,.ADDRTD12 ( ADDRTD12 ) ,.ADDRTD11 ( ADDRTD11 ) ,.ADDRTD10 ( ADDRTD10 )
     ,.ADDRTD9 ( ADDRTD9 ) ,.ADDRTD8 ( ADDRTD8 ) ,.ADDRTD7 ( ADDRTD7 )
     ,.ADDRTD6 ( ADDRTD6 ) ,.ADDRTD5 ( ADDRTD5 ) ,.ADDRTD4 ( ADDRTD4 )
     ,.ADDRTD3 ( ADDRTD3 ) ,.ADDRTD2 ( ADDRTD2 ) ,.ADDRTD1 ( ADDRTD1 )
     ,.ADDRPINRD ( ADDRPINRD ) ,.ADDRPINMD ( ADDRPINMD ) ,.ADDRPINLV ( ADDRPINLV )
     ,.ICEDI0 ( ICEDI0 ) ,.ICEWR ( ICEWR ) ,.PSEUDOON31 ( PSEUDOON31 )
     ,.PSEUDOON23 ( PSEUDOON23 ) ,.PSEUDOON15 ( PSEUDOON15 ) ,.PSEUDOON30 ( PSEUDOON30 )
     ,.PSEUDOON22 ( PSEUDOON22 ) ,.PSEUDOON14 ( PSEUDOON14 ) ,.PSEUDOON29 ( PSEUDOON29 )
     ,.PSEUDOON28 ( PSEUDOON28 ) ,.PSEUDOON27 ( PSEUDOON27 ) ,.PSEUDOON19 ( PSEUDOON19 )
     ,.PSEUDOON26 ( PSEUDOON26 ) ,.PSEUDOON18 ( PSEUDOON18 ) ,.PSEUDOON25 ( PSEUDOON25 )
     ,.PSEUDOON17 ( PSEUDOON17 ) ,.PSEUDOON24 ( PSEUDOON24 ) ,.PSEUDOON16 ( PSEUDOON16 )
     ,.PSEUDOON21 ( PSEUDOON21 ) ,.PSEUDOON13 ( PSEUDOON13 ) ,.PSEUDOON20 ( PSEUDOON20 )
     ,.PSEUDOON12 ( PSEUDOON12 ) ,.PSEUDOON11 ( PSEUDOON11 ) ,.PSEUDOON10 ( PSEUDOON10 )
     ,.PSEUDOON9 ( PSEUDOON9 ) ,.PSEUDOON8 ( PSEUDOON8 ) ,.ICEMSKRETRY ( ICEMSKRETRY )
     ,.ICEMSKTRAP ( ICEMSKTRAP ) ,.ICEMSKWAIT ( ICEMSKWAIT ) ,.IDVER31 ( IDVER31 )
     ,.IDVER23 ( IDVER23 ) ,.IDVER15 ( IDVER15 ) ,.IDVER30 ( IDVER30 )
     ,.IDVER22 ( IDVER22 ) ,.IDVER14 ( IDVER14 ) ,.IDVER29 ( IDVER29 )
     ,.IDVER28 ( IDVER28 ) ,.IDVER27 ( IDVER27 ) ,.IDVER19 ( IDVER19 )
     ,.IDVER26 ( IDVER26 ) ,.IDVER18 ( IDVER18 ) ,.IDVER25 ( IDVER25 )
     ,.IDVER17 ( IDVER17 ) ,.IDVER24 ( IDVER24 ) ,.IDVER16 ( IDVER16 )
     ,.IDVER21 ( IDVER21 ) ,.IDVER13 ( IDVER13 ) ,.IDVER20 ( IDVER20 )
     ,.IDVER12 ( IDVER12 ) ,.IDVER11 ( IDVER11 ) ,.IDVER10 ( IDVER10 )
     ,.IDVER9 ( IDVER9 ) ,.IDVER8 ( IDVER8 ) ,.IDVER7 ( IDVER7 ) ,.IDVER6 ( IDVER6 )
     ,.IDVER5 ( IDVER5 ) ,.IDVER4 ( IDVER4 ) ,.IDVER3 ( IDVER3 ) ,.IDVER2 ( IDVER2 )
     ,.IDVER1 ( IDVER1 ) ,.IDVER0 ( IDVER0 ) ,.EROMPD32 ( EROMPD32 ) ,.EROMPD33 ( EROMPD33 )
     ,.EROMPD34 ( EROMPD34 ) ,.EROMPD35 ( EROMPD35 ) ,.CPURCLK1 ( CPURCLK1 )
     ,.CPURCLK2 ( CPURCLK2 ) ,.SOFTBRK ( SOFTBRK ) ,.OCDMOD ( OCDMOD )
     ,.SBANDOCD ( SBANDOCD ) ,.CLK60MHZLOCK ( CLK60MHZLOCK ) ,.DCER_OUT ( DCER_OUT )
     ,.DDIS_OUT ( DDIS_OUT ) ,.DFCLK_OUT ( DFCLK_OUT ) ,.DMRG00_OUT ( DMRG00_OUT )
     ,.DMRG01_OUT ( DMRG01_OUT ) ,.DMRG10_OUT ( DMRG10_OUT ) ,.DMRG11_OUT ( DMRG11_OUT )
     ,.DMRG12_OUT ( DMRG12_OUT ) ,.DRDCLKP1_OUT ( DRDCLKP1_OUT ) ,.DREAD_OUT ( DREAD_OUT )
     ,.DSER_OUT ( DSER_OUT ) ,.DWWR_OUT ( DWWR_OUT ) ,.LVISEL ( LVISEL )
    
  ) ; 
endmodule

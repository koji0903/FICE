module DriveChangeB_Replace(a);
   input 	   a;
endmodule // DriveChangeB
module ConnectA(I);
   input I;   
endmodule // ConnectA

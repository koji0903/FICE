// created by mkice.pl ver1.0

module chiptop_other (
	ADBIONB ,ADCMP ,ADCPON ,ADINL5V ,ADOFC ,ADPDB ,DSRCUT ,DTRMCP010 ,DTRMCP011 ,DTRMCP012
	,DTRMCP013 ,DTRMCP014 ,HVPPTS1 ,INCDECWS0 ,INCDECWS1 ,MODENOP ,MODERD ,MODEWR ,MUTEST ,PSTN
	,R0A0 ,R0A1 ,R0A2 ,R0A3 ,R0A4 ,R0A5 ,R0FLAGZ ,SELIN1 ,SELTAR ,SRCUTCP
	,TRMCP010 ,TRMCP011 ,TRMCP012 ,TRMCP013 ,TRMCP014 ,TRMRD2 ,TSTN ,VBRESZCP ,VPBIAS ,VPPTS1
	,VREGMV ,VREGRMV ,WDWR
);

	input	ADBIONB ,ADCMP ,ADCPON ,ADINL5V ,ADOFC ,ADPDB ,DSRCUT ,DTRMCP010
		,DTRMCP011 ,DTRMCP012 ,DTRMCP013 ,DTRMCP014 ,HVPPTS1 ,INCDECWS0 ,INCDECWS1 ,MODENOP
		,MODERD ,MODEWR ,MUTEST ,PSTN ,R0A0 ,R0A1 ,R0A2 ,R0A3
		,R0A4 ,R0A5 ,R0FLAGZ ,SELIN1 ,SELTAR ,SRCUTCP ,TRMCP010 ,TRMCP011
		,TRMCP012 ,TRMCP013 ,TRMCP014 ,TRMRD2 ,TSTN ,VBRESZCP ,VPBIAS ,VPPTS1
		,VREGMV ,VREGRMV ,WDWR ;

endmodule


//  file name   ... /proj/78k0r_11/78k0r_kx4/_ice/_make_chip/_1chip_v2.3/_library/d78f1070_cf1.02_eva.hdl
//  top module  ... /proj/78k0r_11/78k0r_kx4/_ice/_make_chip/_1chip_v2.3/_library/d78f1070_cf1.02_eva.hdl D78F1070_EVA
//  version     ... 2.00
//  designer    ... T.Tsunoda
//  refer to    ... make_chip.para

module D78F1070_EVA (
  ADEOCB ,ADSAR0 ,P52DIN ,P60DIN ,ADSAR1 ,P27ENI ,P43ENI ,P51ENI ,ADSAR2 ,ADSAR3 ,ADSAR4
 ,ADSAR5 ,ADSAR6 ,ADSAR7 ,P27ENO ,P43ENO ,P51ENO ,ADSAR8 ,P53DIN ,P61DIN ,ADSAR9
 ,P52ENI ,P60ENI ,DRO00 ,DRO01 ,DRO010 ,DRO011 ,DRO02 ,DRO03 ,DRO04 ,FIHFL
 ,DRO05 ,DRO06 ,DRO07 ,DRO08 ,DRO09 ,EIRAMO0 ,EIRAMO1 ,FIHOCD ,HVIN ,LVIOUTZNF
 ,MDRRAM0 ,MDRRAM1 ,MDRRAM10 ,MDRRAM11 ,MDRRAM12 ,MDRRAM13 ,MDRRAM14 ,MDRRAM15 ,MDRRAM2 ,MDRRAM3
 ,MDRRAM4 ,MDRRAM5 ,MDRRAM6 ,FRQSEL0 ,MDRRAM7 ,FRQSEL1 ,MDRRAM8 ,FRQSEL2 ,MDRRAM9 ,FRQSEL3
 ,MODE0 ,MODE1 ,OSCOUTM ,OSCOUTS ,P00DIN ,P01DIN ,P02DIN ,P10DIN ,P03DIN ,P11DIN
 ,P04DIN ,P12DIN ,P20DIN ,P05DIN ,P13DIN ,P21DIN ,P06DIN ,P14DIN ,P22DIN ,P30DIN
 ,P120DIN ,P137DIN ,P140DIN ,P141DIN ,P146DIN ,P147DIN ,P147SELIN1B5V ,P15DIN ,P23DIN ,P31DIN
 ,P16DIN ,P24DIN ,P40DIN ,P17DIN ,P25DIN ,P41DIN ,P26DIN ,P42DIN ,P50DIN ,P27DIN
 ,P43DIN ,P51DIN ,P40SELIN1B5V ,P54DIN ,P62DIN ,P70DIN ,DGEN00 ,P55DIN ,P63DIN ,P71DIN
 ,P72DIN ,P73DIN ,P74DIN ,P75DIN ,P76DIN ,P77DIN ,POCREL ,RESETB ,POCREL5V ,POCRELNF
 ,R15KOUT ,R32MOUT ,RESETINBNF ,RO00 ,PID0 ,MDW6 ,RO01 ,PID1 ,MDW7 ,RO010
 ,PID10 ,RO011 ,PID11 ,RO012 ,RO020 ,PID20 ,PID12 ,CPURD ,RO013 ,RO021
 ,PID21 ,PID13 ,RO014 ,RO022 ,RO030 ,PID30 ,PID22 ,PID14 ,RO110 ,RO015
 ,RO023 ,RO031 ,PID31 ,PID23 ,PID15 ,RO111 ,RO016 ,RO024 ,RO032 ,PID24
 ,PID16 ,RO120 ,RO112 ,RO017 ,RO025 ,RO033 ,PID25 ,PID17 ,RO121 ,RO113
 ,RO018 ,RO026 ,RO034 ,PID26 ,PID18 ,RO130 ,RO122 ,RO114 ,RO019 ,RO027
 ,RO035 ,PID27 ,PID19 ,RO131 ,RO123 ,RO115 ,RO02 ,PID2 ,RO10 ,MDW8
 ,RO028 ,RO036 ,PID28 ,RO132 ,RO124 ,RO116 ,RO029 ,RO037 ,PID29 ,RO133
 ,RO125 ,RO117 ,RO03 ,PID3 ,RO11 ,MDW9 ,RO04 ,PID4 ,RO12 ,RO05
 ,PID5 ,RO13 ,RO06 ,PID6 ,RO14 ,RO07 ,PID7 ,RO15 ,RO08 ,PID8
 ,RO16 ,RO09 ,PID9 ,RO17 ,RPERR ,RTCCLK ,STN ,TRESET ,VREG ,X1DIN
 ,RO136 ,RO128 ,EXMA2 ,X2DIN ,XT1DIN ,XT2DIN ,A10 ,A11 ,A12 ,A13
 ,A14 ,A15 ,A2 ,A3 ,A4 ,A5 ,A6 ,A7 ,A8 ,A9
 ,ADBIONB ,ADCHSEL0 ,ADCHSEL1 ,ADCHSEL2 ,ADCHSEL3 ,ADCHSEL4 ,ADCLK ,ADCMP ,ADCPON ,ADGSELMOD
 ,ADINL5V ,ADOFC ,ADPDB ,ADS1 ,ADTESMOD0 ,ADTESMOD1 ,ADTESMOD2 ,ADVSELMOD0 ,ADVSELMOD1 ,AMPH
 ,PC16 ,AMPHS0 ,AMPHS1 ,AMPSEL ,BEU0 ,MA10 ,BEU1 ,MA11 ,BEU2 ,MA12
 ,BFA ,BG1ST ,BG2ADEN ,BG2ADSEL ,BGRT0 ,BGRT1 ,BGRT10 ,BGRT2 ,BGRT3 ,BGRT4
 ,BGRT5 ,BGRT6 ,BGRT7 ,BGRT8 ,BGRT9 ,BRSAM ,CPUCLKEN ,CTRIM0 ,CTRIM1 ,CTRIM2
 ,CTRIM3 ,CTRIM4 ,CTRIM5 ,CTRIM6 ,DA0 ,AF2 ,DA1 ,AF3 ,DA10 ,AF14
 ,DA11 ,AF15 ,DA2 ,AF4 ,DA3 ,AF5 ,DA4 ,CE0 ,AF6 ,DA5
 ,CE1 ,AF7 ,DA6 ,AF8 ,DA7 ,AF9 ,DA8 ,DA9 ,DSRCUT ,DTRMCP010
 ,DTRMCP011 ,DTRMCP012 ,DTRMCP013 ,DTRMCP014 ,DW0 ,MA8 ,DW1 ,MA9 ,DW10 ,DW11
 ,DW12 ,DW20 ,DW13 ,DW21 ,ALT1 ,DW14 ,DW22 ,DW30 ,DW15 ,DW23
 ,DW31 ,DW16 ,DW24 ,DW32 ,DW17 ,DW25 ,DW33 ,DDIS ,DW18 ,DW26
 ,DW34 ,PA10 ,DW19 ,DW27 ,DW35 ,PA11 ,DW2 ,DW28 ,DW36 ,PA12
 ,DW29 ,DW37 ,PA13 ,DW3 ,DW4 ,DW5 ,DW6 ,PA2 ,DW7 ,PA3
 ,DIS ,DW8 ,PA4 ,PC0 ,DW9 ,PA5 ,PC1 ,EXA ,EXCLK ,EXCLKS
 ,FCLK2 ,FRSEL0 ,FRSEL1 ,FRSEL2 ,FRSEL3 ,FRSEL4 ,FTRIM0 ,FTRIM1 ,FTRIM2 ,FTRIM3
 ,FTRIM4 ,FTRIM5 ,HVPPTS1 ,INCDECWS0 ,INCDECWS1 ,LOSCTEST ,LVIEN ,LVIS2 ,LVIS0 ,LVIS1
 ,LVIS3 ,LVITEST ,LVITSEL ,MDLYCUT ,MODENOP ,MODERD ,MODEWR ,MSTOP ,MUTEST ,OREGSTP
 ,OSCSEL ,PREFIX ,OSCSELS ,P00DOUT ,P00ENI ,P00ENO ,P00PUON ,P01DOUT ,P01ENI ,P01ENO
 ,P01PUON ,P01SELIN ,P02DOUT ,P10DOUT ,P02ENI ,P10ENI ,P02ENO ,P10ENO ,P02PUON ,P10PUON
 ,P03DOUT ,P11DOUT ,P03ENI ,P11ENI ,P03ENO ,P11ENO ,P03PUON ,P11PUON ,P03SELIN ,P11SELIN
 ,P04DOUT ,P12DOUT ,P20DOUT ,P04ENI ,P12ENI ,P20ENI ,P04ENO ,P12ENO ,P20ENO ,P04PUON
 ,P12PUON ,P04SELIN ,P05DOUT ,P13DOUT ,P21DOUT ,P05ENI ,P13ENI ,P21ENI ,P05ENO ,P13ENO
 ,P21ENO ,P05PUON ,P13PUON ,P06DOUT ,P14DOUT ,P22DOUT ,P30DOUT ,P06ENI ,P14ENI ,P22ENI
 ,P30ENI ,P06ENO ,P14ENO ,P22ENO ,P30ENO ,P06PUON ,P14PUON ,P30PUON ,P10SELIN ,P120DOUT
 ,P120ENI ,P120ENO ,P120PUON ,P130DOUT ,P130ENO ,P137ENI ,P13SELIN ,P140DOUT ,P140ENI ,P140ENO
 ,P140PUON ,P141DOUT ,P141ENI ,P141ENO ,P141PUON ,P146DOUT ,P146ENI ,P146ENO ,P146PUON ,P147DOUT
 ,P147ENI ,P147ENO ,P147PUON ,P14SELIN ,P15DOUT ,P23DOUT ,P31DOUT ,P15ENI ,P23ENI ,P31ENI
 ,P15ENO ,P23ENO ,P31ENO ,P15PUON ,P31PUON ,P15SELIN ,P16DOUT ,P24DOUT ,P40DOUT ,P16ENI
 ,P24ENI ,P40ENI ,P16ENO ,P24ENO ,P40ENO ,P16PUON ,P40PUON ,P16SELIN ,P17DOUT ,P25DOUT
 ,P41DOUT ,P17ENI ,P25ENI ,P41ENI ,P17ENO ,P25ENO ,P41ENO ,P17PUON ,P41PUON ,P17SELIN
 ,P26DOUT ,P42DOUT ,P50DOUT ,P26ENI ,P42ENI ,P50ENI ,P26ENO ,P42ENO ,P50ENO ,P27DOUT
 ,P43DOUT ,P51DOUT ,P42PUON ,P50PUON ,P43PUON ,P51PUON ,P52DOUT ,P60DOUT ,P52ENO ,P60ENO
 ,P52PUON ,P53DOUT ,P61DOUT ,P53ENI ,P61ENI ,DGEN01 ,P53ENO ,P61ENO ,DGEN07 ,P53PUON
 ,P54DOUT ,P62DOUT ,P70DOUT ,P54ENI ,P62ENI ,P70ENI ,P54ENO ,P62ENO ,P70ENO ,P54PUON
 ,P70PUON ,P55DOUT ,P63DOUT ,P71DOUT ,P55ENI ,P63ENI ,P71ENI ,P55ENO ,P63ENO ,P71ENO
 ,P55PUON ,P71PUON ,P55SELIN ,P72DOUT ,P72ENI ,P72ENO ,P72PUON ,P73DOUT ,P73ENI ,P73ENO
 ,P73PUON ,IDADR24 ,IDADR16 ,P74DOUT ,P74ENI ,P74ENO ,P74PUON ,ICEDO20 ,ICEDO12 ,P75DOUT
 ,P75ENI ,P75ENO ,P75PUON ,P76DOUT ,P76ENI ,P76ENO ,P76PUON ,P77DOUT ,P77ENI ,P77ENO
 ,P77PUON ,PAENB ,PSTN ,R0A0 ,MA14 ,R0A1 ,MA15 ,R0A2 ,R0A3 ,R0A4
 ,R0A5 ,R0FLAGZ ,REG125ST ,REGLC ,REGLV ,RTCCLKEN ,RTRIM0 ,RTRIM1 ,RTRIM2 ,RTRIM3
 ,RTRIM4 ,RTRIM5 ,SELIN1 ,SELTAR ,SRCUTCP ,STOPZ ,TRMCP010 ,TRMCP011 ,TRMCP012 ,TRMCP013
 ,TRMCP014 ,TRMRD2 ,TSTN ,VBRESZCP ,VPBIAS ,XT2ENI ,VPPTS1 ,VREGMV ,VREGRMV ,WDWR
 ,WTRIM0 ,WTRIM1 ,WTRIM2 ,X1ENI ,X2ENI ,XT1ENI ,XTSTOP ,XTWKUP ,reg_adtyp ,A19
 ,A18 ,A17 ,A16 ,SELRO1 ,CLKSEL1 ,ICETMSPMD ,ICETMBTSEL ,RO137 ,RO129 ,EXMA3
 ,FLSPM ,RO135 ,RO127 ,RO119 ,EXMA1 ,RO134 ,RO126 ,RO118 ,EXMA0 ,RO19
 ,RO18 ,DCE0 ,DCLKSEL1 ,DRDCLKC1 ,DA13 ,AF17 ,DA12 ,AF16 ,SLFLASH ,WAITFL2
 ,SVI ,SVVCOUT7 ,SVVCOUT6 ,SVVCOUT5 ,SVVCOUT4 ,SVVCOUT3 ,SVVCOUT2 ,SVVCOUT1 ,SVVCOUT0 ,SVINTACK
 ,SOFTBRK ,ICEMSKNMI ,ICEMSKDBG ,STAGEADR1 ,STAGEADR0 ,SKIPEXE ,PCWAITF ,CPUMASK ,CPUPID1 ,CPUMISAL
 ,FLREAD ,IMDR10 ,FLREADB3 ,FLREADB2 ,FLREADB1 ,FLREADB0 ,FCHRAM ,SLMEM ,SLEXM ,SLBMEM
 ,SPDEC ,SPINC ,SPREL ,IDPOP ,MDW10 ,IMDR2 ,CPUWR ,WDOP ,ICEWAITMEM ,DMAACK
 ,HLTST ,STPST ,INTACK ,OCDWAIT ,SVMOD ,SVMODF ,DRDCLK ,SLDFLASH ,ICECSGREGU ,ICEIFA4
 ,ICEIFA3 ,ICEIFA2 ,ICEDO31 ,ICEDO23 ,ICEDO15 ,ICEDO30 ,ICEDO22 ,ICEDO14 ,ICEDO29 ,ICEDO28
 ,ICEDO27 ,ICEDO19 ,ICEDO26 ,ICEDO18 ,ICEDO25 ,ICEDO17 ,ICEDO24 ,ICEDO16 ,ICEDO21 ,ICEDO13
 ,ICEDO11 ,ICEDO10 ,ICEDO9 ,ICEDO8 ,ICEDO7 ,ICEDO6 ,ICEDO5 ,ICEDO4 ,ICEDO3 ,ICEDO2
 ,ICEDO1 ,ICEDO0 ,PA19 ,PC11 ,PA18 ,PC10 ,PA17 ,PA16 ,PA15 ,PA14
 ,PA9 ,PC5 ,PA8 ,PC4 ,PA7 ,PC3 ,PA6 ,PC2 ,PC19 ,PC18
 ,PC17 ,PC15 ,PC14 ,PC13 ,PC12 ,PC9 ,PC8 ,PC7 ,PC6 ,IDADR31
 ,IDADR23 ,IDADR15 ,IDADR30 ,IDADR22 ,IDADR14 ,IDADR29 ,IDADR28 ,IDADR27 ,IDADR19 ,IDADR26
 ,IDADR18 ,IDADR25 ,IDADR17 ,IDADR21 ,IDADR13 ,IDADR20 ,IDADR12 ,IDADR11 ,IDADR10 ,IDADR9
 ,IDADR8 ,IDADR7 ,IDADR6 ,IDADR5 ,IDADR4 ,IDADR3 ,IDADR2 ,IDADR1 ,IDADR0 ,MA13
 ,MA7 ,MA6 ,MA5 ,MA4 ,MA3 ,MA2 ,CER ,MA1 ,MA0 ,MDW15
 ,IMDR7 ,MDW14 ,IMDR6 ,MDW13 ,IMDR5 ,MDW12 ,IMDR4 ,MDW11 ,IMDR3 ,MDW5
 ,MDW4 ,MDW3 ,MDW2 ,MDW1 ,MDW0 ,EXCH ,IMDR15 ,IMDR14 ,IMDR13 ,IMDR12
 ,IMDR11 ,IMDR9 ,IMDR8 ,IMDR1 ,IMDR0 ,CPUPID31 ,CPUPID23 ,CPUPID15 ,CPUPID30 ,CPUPID22
 ,CPUPID14 ,CPUPID29 ,CPUPID28 ,CPUPID27 ,CPUPID19 ,CPUPID26 ,CPUPID18 ,CPUPID25 ,CPUPID17 ,CPUPID24
 ,CPUPID16 ,CPUPID21 ,CPUPID13 ,CPUPID20 ,CPUPID12 ,CPUPID11 ,CPUPID10 ,CPUPID9 ,CPUPID8 ,CPUPID7
 ,CPUPID6 ,CPUPID5 ,CPUPID4 ,CPUPID3 ,CPUPID2 ,CPUPID0 ,FLSIZE3 ,FLSIZE2 ,FLSIZE1 ,FLSIZE0
 ,RAMSIZE7 ,RAMSIZE6 ,RAMSIZE5 ,RAMSIZE4 ,RAMSIZE3 ,RAMSIZE2 ,RAMSIZE1 ,RAMSIZE0 ,BFSIZE3 ,BFSIZE2
 ,BFSIZE1 ,BFSIZE0 ,BMSIZE3 ,BMSIZE2 ,BMSIZE1 ,BMSIZE0 ,DFSIZE1 ,DFSIZE0 ,ICEMKLVI ,ICEMKWDT
 ,ICEMKSRQ ,RESB ,FCLKRT ,CIBRESRQ ,CIBRESRQICE ,FCLK1 ,TMSPMD ,TMBTSEL ,BTFLG ,READ
 ,RDCLKP1 ,SER ,WED ,WWR ,MRG00 ,MRG01 ,MRG10 ,MRG11 ,MRG12 ,PROGI
 ,ICEFLERR ,ICENOECC ,DCER ,DSER ,DWWR ,DWED ,DMRG00 ,DMRG01 ,DMRG10 ,DMRG11
 ,DMRG12 ,DREAD ,AF19 ,AF18 ,AF13 ,AF12 ,AF11 ,AF10 ,AF1 ,AF0
 ,OCDMOD ,ICECK60M ,CLK60MHZ ,CLK60M ,GDRAMWR ,IAWRES ,SVSTOPIAW ,CPUWRIAW ,PSEUDOON10 ,PSEUDOON1
 ,SVSTOPICE ,SVSTOP ,SVPERI0ICE ,SVPERI0 ,SVPERI1ICE ,SVPERI1 ,MONMD ,MONSVMOD ,STBRELE ,STBRELEICE
 ,FRQSEL4 ,R32MSTP ,REQOCD ,REQFL ,TSELOREG ,TSELIRES ,TTEMP ,R15KSTPZ ,SYSRESB ,OPLVIMDS1
 ,OPLVIMDS0 ,SCANCLKICE ,SCANMODEICE ,SCANRESZICE ,SCANENICE ,SCANCLK ,SCANMODE ,SCANRESZ ,SCANEN ,CKSMER
 ,ICEDATAFLT ,ICEDMAFLT ,ICEFETCHFLT ,ICESVSTOP ,TIIDER ,PSEUDOTIIDER ,ICECKSMER ,CSPDTFLP ,CSPDTFLG ,RAMSIZE7ICE
 ,RAMSIZE6ICE ,RAMSIZE5ICE ,RAMSIZE4ICE ,RAMSIZE3ICE ,RAMSIZE2ICE ,RAMSIZE1ICE ,RAMSIZE0ICE ,FLSIZE3ICE ,FLSIZE2ICE ,FLSIZE1ICE
 ,FLSIZE0ICE ,DFSIZE1ICE ,DFSIZE0ICE ,SYSRSOUTB ,PIO00 ,PIO01 ,PIO02 ,PIO10 ,PIO03 ,PIO11
 ,PIO04 ,PIO12 ,PIO20 ,PIO05 ,PIO13 ,PIO21 ,PIO06 ,PIO14 ,PIO22 ,PIO30
 ,PIO15 ,PIO23 ,PIO31 ,PIO16 ,PIO24 ,PIO40 ,PIO17 ,PIO25 ,PIO41 ,PIO26
 ,PIO42 ,PIO50 ,PIO27 ,PIO43 ,PIO51 ,PIO52 ,PIO60 ,PIO53 ,PIO61 ,PIO54
 ,PIO62 ,PIO70 ,PIO55 ,PIO63 ,PIO71 ,PIO72 ,PIO73 ,PIO74 ,PIO75 ,PIO76
 ,PIO77 ,PIO120 ,PIO121 ,PIO122 ,PIO130 ,PIO123 ,PIO124 ,PIO140 ,PIO137 ,PIO141
 ,PIO146 ,PIO147 ,PRESADCZ ,DGEN06 ,DGEN05 ,DGEN04 ,DGEN03 ,DGEN02
);

  input ADEOCB ;
  input ADSAR0 ;
  input P52DIN ;
  input P60DIN ;
  input ADSAR1 ;
  input ADSAR2 ;
  input ADSAR3 ;
  input ADSAR4 ;
  input ADSAR5 ;
  input ADSAR6 ;
  input ADSAR7 ;
  input ADSAR8 ;
  input P53DIN ;
  input P61DIN ;
  input ADSAR9 ;
  input DRO00 ;
  input DRO01 ;
  input DRO010 ;
  input DRO011 ;
  input DRO02 ;
  input DRO03 ;
  input DRO04 ;
  input FIHFL ;
  input DRO05 ;
  input DRO06 ;
  input DRO07 ;
  input DRO08 ;
  input DRO09 ;
  input EIRAMO0 ;
  input EIRAMO1 ;
  input FIHOCD ;
  input HVIN ;
  input LVIOUTZNF ;
  input MDRRAM0 ;
  input MDRRAM1 ;
  input MDRRAM10 ;
  input MDRRAM11 ;
  input MDRRAM12 ;
  input MDRRAM13 ;
  input MDRRAM14 ;
  input MDRRAM15 ;
  input MDRRAM2 ;
  input MDRRAM3 ;
  input MDRRAM4 ;
  input MDRRAM5 ;
  input MDRRAM6 ;
  input MDRRAM7 ;
  input MDRRAM8 ;
  input MDRRAM9 ;
  input MODE0 ;
  input MODE1 ;
  input OSCOUTM ;
  input OSCOUTS ;
  input P00DIN ;
  input P01DIN ;
  input P02DIN ;
  input P10DIN ;
  input P03DIN ;
  input P11DIN ;
  input P04DIN ;
  input P12DIN ;
  input P20DIN ;
  input P05DIN ;
  input P13DIN ;
  input P21DIN ;
  input P06DIN ;
  input P14DIN ;
  input P22DIN ;
  input P30DIN ;
  input P120DIN ;
  input P137DIN ;
  input P140DIN ;
  input P141DIN ;
  input P146DIN ;
  input P147DIN ;
  input P147SELIN1B5V ;
  input P15DIN ;
  input P23DIN ;
  input P31DIN ;
  input P16DIN ;
  input P24DIN ;
  input P40DIN ;
  input P17DIN ;
  input P25DIN ;
  input P41DIN ;
  input P26DIN ;
  input P42DIN ;
  input P50DIN ;
  input P27DIN ;
  input P43DIN ;
  input P51DIN ;
  input P40SELIN1B5V ;
  input P54DIN ;
  input P62DIN ;
  input P70DIN ;
  input P55DIN ;
  input P63DIN ;
  input P71DIN ;
  input P72DIN ;
  input P73DIN ;
  input P74DIN ;
  input P75DIN ;
  input P76DIN ;
  input P77DIN ;
  input POCREL ;
  input POCREL5V ;
  input POCRELNF ;
  input R15KOUT ;
  input R32MOUT ;
  input RESETINBNF ;
  input RO00 ;
  input RO01 ;
  input RO010 ;
  input RO011 ;
  input RO012 ;
  input RO020 ;
  input RO013 ;
  input RO021 ;
  input RO014 ;
  input RO022 ;
  input RO030 ;
  input RO110 ;
  input RO015 ;
  input RO023 ;
  input RO031 ;
  input RO111 ;
  input RO016 ;
  input RO024 ;
  input RO032 ;
  input RO120 ;
  input RO112 ;
  input RO017 ;
  input RO025 ;
  input RO033 ;
  input RO121 ;
  input RO113 ;
  input RO018 ;
  input RO026 ;
  input RO034 ;
  input RO130 ;
  input RO122 ;
  input RO114 ;
  input RO019 ;
  input RO027 ;
  input RO035 ;
  input RO131 ;
  input RO123 ;
  input RO115 ;
  input RO02 ;
  input RO10 ;
  input RO028 ;
  input RO036 ;
  input RO132 ;
  input RO124 ;
  input RO116 ;
  input RO029 ;
  input RO037 ;
  input RO133 ;
  input RO125 ;
  input RO117 ;
  input RO03 ;
  input RO11 ;
  input RO04 ;
  input RO12 ;
  input RO05 ;
  input RO13 ;
  input RO06 ;
  input RO14 ;
  input RO07 ;
  input RO15 ;
  input RO08 ;
  input RO16 ;
  input RO09 ;
  input RO17 ;
  input RPERR ;
  input RTCCLK ;
  input STN ;
  input TRESET ;
  input VREG ;
  input X1DIN ;
  input RO136 ;
  input RO128 ;
  input X2DIN ;
  input XT1DIN ;
  input XT2DIN ;
  input ICETMSPMD ;
  input ICETMBTSEL ;
  input RO137 ;
  input RO129 ;
  input RO135 ;
  input RO127 ;
  input RO119 ;
  input RO134 ;
  input RO126 ;
  input RO118 ;
  input RO19 ;
  input RO18 ;
  input WAITFL2 ;
  input SVI ;
  input SVVCOUT7 ;
  input SVVCOUT6 ;
  input SVVCOUT5 ;
  input SVVCOUT4 ;
  input SVVCOUT3 ;
  input SVVCOUT2 ;
  input SVVCOUT1 ;
  input SVVCOUT0 ;
  input ICEMSKNMI ;
  input ICEMSKDBG ;
  input CPUPID1 ;
  input ICEWAITMEM ;
  input ICECSGREGU ;
  input ICEIFA4 ;
  input ICEIFA3 ;
  input ICEIFA2 ;
  input CPUPID31 ;
  input CPUPID23 ;
  input CPUPID15 ;
  input CPUPID30 ;
  input CPUPID22 ;
  input CPUPID14 ;
  input CPUPID29 ;
  input CPUPID28 ;
  input CPUPID27 ;
  input CPUPID19 ;
  input CPUPID26 ;
  input CPUPID18 ;
  input CPUPID25 ;
  input CPUPID17 ;
  input CPUPID24 ;
  input CPUPID16 ;
  input CPUPID21 ;
  input CPUPID13 ;
  input CPUPID20 ;
  input CPUPID12 ;
  input CPUPID11 ;
  input CPUPID10 ;
  input CPUPID9 ;
  input CPUPID8 ;
  input CPUPID7 ;
  input CPUPID6 ;
  input CPUPID5 ;
  input CPUPID4 ;
  input CPUPID3 ;
  input CPUPID2 ;
  input CPUPID0 ;
  input FLSIZE3 ;
  input FLSIZE2 ;
  input FLSIZE1 ;
  input FLSIZE0 ;
  input RAMSIZE7 ;
  input RAMSIZE6 ;
  input RAMSIZE5 ;
  input RAMSIZE4 ;
  input RAMSIZE3 ;
  input RAMSIZE2 ;
  input RAMSIZE1 ;
  input RAMSIZE0 ;
  input BFSIZE3 ;
  input BFSIZE2 ;
  input BFSIZE1 ;
  input BFSIZE0 ;
  input BMSIZE3 ;
  input BMSIZE2 ;
  input BMSIZE1 ;
  input BMSIZE0 ;
  input DFSIZE1 ;
  input DFSIZE0 ;
  input ICEMKLVI ;
  input ICEMKWDT ;
  input ICEMKSRQ ;
  input CIBRESRQICE ;
  input ICEFLERR ;
  input ICENOECC ;
  input ICECK60M ;
  input CLK60MHZ ;
  input CLK60M ;
  input SVSTOPIAW ;
  input CPUWRIAW ;
  input PSEUDOON10 ;
  input PSEUDOON1 ;
  input SVSTOP ;
  input SVPERI0 ;
  input SVPERI1 ;
  input MONSVMOD ;
  input STBRELEICE ;
  input SCANCLK ;
  input SCANMODE ;
  input SCANRESZ ;
  input SCANEN ;
  input ICEDATAFLT ;
  input ICEDMAFLT ;
  input ICEFETCHFLT ;
  input ICESVSTOP ;
  input PSEUDOTIIDER ;
  input ICECKSMER ;
  input CSPDTFLG ;
  input SYSRSOUTB ;

  output P27ENI ;
  output P43ENI ;
  output P51ENI ;
  output P27ENO ;
  output P43ENO ;
  output P51ENO ;
  output P52ENI ;
  output P60ENI ;
  output FRQSEL0 ;
  output FRQSEL1 ;
  output FRQSEL2 ;
  output FRQSEL3 ;
  output DGEN00 ;
  output RESETB ;
  output PID0 ;
  output MDW6 ;
  output PID1 ;
  output MDW7 ;
  output PID10 ;
  output PID11 ;
  output PID20 ;
  output PID12 ;
  output CPURD ;
  output PID21 ;
  output PID13 ;
  output PID30 ;
  output PID22 ;
  output PID14 ;
  output PID31 ;
  output PID23 ;
  output PID15 ;
  output PID24 ;
  output PID16 ;
  output PID25 ;
  output PID17 ;
  output PID26 ;
  output PID18 ;
  output PID27 ;
  output PID19 ;
  output PID2 ;
  output MDW8 ;
  output PID28 ;
  output PID29 ;
  output PID3 ;
  output MDW9 ;
  output PID4 ;
  output PID5 ;
  output PID6 ;
  output PID7 ;
  output PID8 ;
  output PID9 ;
  output EXMA2 ;
  output A10 ;
  output A11 ;
  output A12 ;
  output A13 ;
  output A14 ;
  output A15 ;
  output A2 ;
  output A3 ;
  output A4 ;
  output A5 ;
  output A6 ;
  output A7 ;
  output A8 ;
  output A9 ;
  output ADBIONB ;
  output ADCHSEL0 ;
  output ADCHSEL1 ;
  output ADCHSEL2 ;
  output ADCHSEL3 ;
  output ADCHSEL4 ;
  output ADCLK ;
  output ADCMP ;
  output ADCPON ;
  output ADGSELMOD ;
  output ADINL5V ;
  output ADOFC ;
  output ADPDB ;
  output ADS1 ;
  output ADTESMOD0 ;
  output ADTESMOD1 ;
  output ADTESMOD2 ;
  output ADVSELMOD0 ;
  output ADVSELMOD1 ;
  output AMPH ;
  output PC16 ;
  output AMPHS0 ;
  output AMPHS1 ;
  output AMPSEL ;
  output BEU0 ;
  output MA10 ;
  output BEU1 ;
  output MA11 ;
  output BEU2 ;
  output MA12 ;
  output BFA ;
  output BG1ST ;
  output BG2ADEN ;
  output BG2ADSEL ;
  output BGRT0 ;
  output BGRT1 ;
  output BGRT10 ;
  output BGRT2 ;
  output BGRT3 ;
  output BGRT4 ;
  output BGRT5 ;
  output BGRT6 ;
  output BGRT7 ;
  output BGRT8 ;
  output BGRT9 ;
  output BRSAM ;
  output CPUCLKEN ;
  output CTRIM0 ;
  output CTRIM1 ;
  output CTRIM2 ;
  output CTRIM3 ;
  output CTRIM4 ;
  output CTRIM5 ;
  output CTRIM6 ;
  output DA0 ;
  output AF2 ;
  output DA1 ;
  output AF3 ;
  output DA10 ;
  output AF14 ;
  output DA11 ;
  output AF15 ;
  output DA2 ;
  output AF4 ;
  output DA3 ;
  output AF5 ;
  output DA4 ;
  output CE0 ;
  output AF6 ;
  output DA5 ;
  output CE1 ;
  output AF7 ;
  output DA6 ;
  output AF8 ;
  output DA7 ;
  output AF9 ;
  output DA8 ;
  output DA9 ;
  output DSRCUT ;
  output DTRMCP010 ;
  output DTRMCP011 ;
  output DTRMCP012 ;
  output DTRMCP013 ;
  output DTRMCP014 ;
  output DW0 ;
  output MA8 ;
  output DW1 ;
  output MA9 ;
  output DW10 ;
  output DW11 ;
  output DW12 ;
  output DW20 ;
  output DW13 ;
  output DW21 ;
  output ALT1 ;
  output DW14 ;
  output DW22 ;
  output DW30 ;
  output DW15 ;
  output DW23 ;
  output DW31 ;
  output DW16 ;
  output DW24 ;
  output DW32 ;
  output DW17 ;
  output DW25 ;
  output DW33 ;
  output DDIS ;
  output DW18 ;
  output DW26 ;
  output DW34 ;
  output PA10 ;
  output DW19 ;
  output DW27 ;
  output DW35 ;
  output PA11 ;
  output DW2 ;
  output DW28 ;
  output DW36 ;
  output PA12 ;
  output DW29 ;
  output DW37 ;
  output PA13 ;
  output DW3 ;
  output DW4 ;
  output DW5 ;
  output DW6 ;
  output PA2 ;
  output DW7 ;
  output PA3 ;
  output DIS ;
  output DW8 ;
  output PA4 ;
  output PC0 ;
  output DW9 ;
  output PA5 ;
  output PC1 ;
  output EXA ;
  output EXCLK ;
  output EXCLKS ;
  output FCLK2 ;
  output FRSEL0 ;
  output FRSEL1 ;
  output FRSEL2 ;
  output FRSEL3 ;
  output FRSEL4 ;
  output FTRIM0 ;
  output FTRIM1 ;
  output FTRIM2 ;
  output FTRIM3 ;
  output FTRIM4 ;
  output FTRIM5 ;
  output HVPPTS1 ;
  output INCDECWS0 ;
  output INCDECWS1 ;
  output LOSCTEST ;
  output LVIEN ;
  output LVIS2 ;
  output LVIS0 ;
  output LVIS1 ;
  output LVIS3 ;
  output LVITEST ;
  output LVITSEL ;
  output MDLYCUT ;
  output MODENOP ;
  output MODERD ;
  output MODEWR ;
  output MSTOP ;
  output MUTEST ;
  output OREGSTP ;
  output OSCSEL ;
  output PREFIX ;
  output OSCSELS ;
  output P00DOUT ;
  output P00ENI ;
  output P00ENO ;
  output P00PUON ;
  output P01DOUT ;
  output P01ENI ;
  output P01ENO ;
  output P01PUON ;
  output P01SELIN ;
  output P02DOUT ;
  output P10DOUT ;
  output P02ENI ;
  output P10ENI ;
  output P02ENO ;
  output P10ENO ;
  output P02PUON ;
  output P10PUON ;
  output P03DOUT ;
  output P11DOUT ;
  output P03ENI ;
  output P11ENI ;
  output P03ENO ;
  output P11ENO ;
  output P03PUON ;
  output P11PUON ;
  output P03SELIN ;
  output P11SELIN ;
  output P04DOUT ;
  output P12DOUT ;
  output P20DOUT ;
  output P04ENI ;
  output P12ENI ;
  output P20ENI ;
  output P04ENO ;
  output P12ENO ;
  output P20ENO ;
  output P04PUON ;
  output P12PUON ;
  output P04SELIN ;
  output P05DOUT ;
  output P13DOUT ;
  output P21DOUT ;
  output P05ENI ;
  output P13ENI ;
  output P21ENI ;
  output P05ENO ;
  output P13ENO ;
  output P21ENO ;
  output P05PUON ;
  output P13PUON ;
  output P06DOUT ;
  output P14DOUT ;
  output P22DOUT ;
  output P30DOUT ;
  output P06ENI ;
  output P14ENI ;
  output P22ENI ;
  output P30ENI ;
  output P06ENO ;
  output P14ENO ;
  output P22ENO ;
  output P30ENO ;
  output P06PUON ;
  output P14PUON ;
  output P30PUON ;
  output P10SELIN ;
  output P120DOUT ;
  output P120ENI ;
  output P120ENO ;
  output P120PUON ;
  output P130DOUT ;
  output P130ENO ;
  output P137ENI ;
  output P13SELIN ;
  output P140DOUT ;
  output P140ENI ;
  output P140ENO ;
  output P140PUON ;
  output P141DOUT ;
  output P141ENI ;
  output P141ENO ;
  output P141PUON ;
  output P146DOUT ;
  output P146ENI ;
  output P146ENO ;
  output P146PUON ;
  output P147DOUT ;
  output P147ENI ;
  output P147ENO ;
  output P147PUON ;
  output P14SELIN ;
  output P15DOUT ;
  output P23DOUT ;
  output P31DOUT ;
  output P15ENI ;
  output P23ENI ;
  output P31ENI ;
  output P15ENO ;
  output P23ENO ;
  output P31ENO ;
  output P15PUON ;
  output P31PUON ;
  output P15SELIN ;
  output P16DOUT ;
  output P24DOUT ;
  output P40DOUT ;
  output P16ENI ;
  output P24ENI ;
  output P40ENI ;
  output P16ENO ;
  output P24ENO ;
  output P40ENO ;
  output P16PUON ;
  output P40PUON ;
  output P16SELIN ;
  output P17DOUT ;
  output P25DOUT ;
  output P41DOUT ;
  output P17ENI ;
  output P25ENI ;
  output P41ENI ;
  output P17ENO ;
  output P25ENO ;
  output P41ENO ;
  output P17PUON ;
  output P41PUON ;
  output P17SELIN ;
  output P26DOUT ;
  output P42DOUT ;
  output P50DOUT ;
  output P26ENI ;
  output P42ENI ;
  output P50ENI ;
  output P26ENO ;
  output P42ENO ;
  output P50ENO ;
  output P27DOUT ;
  output P43DOUT ;
  output P51DOUT ;
  output P42PUON ;
  output P50PUON ;
  output P43PUON ;
  output P51PUON ;
  output P52DOUT ;
  output P60DOUT ;
  output P52ENO ;
  output P60ENO ;
  output P52PUON ;
  output P53DOUT ;
  output P61DOUT ;
  output P53ENI ;
  output P61ENI ;
  output DGEN01 ;
  output P53ENO ;
  output P61ENO ;
  output DGEN07 ;
  output P53PUON ;
  output P54DOUT ;
  output P62DOUT ;
  output P70DOUT ;
  output P54ENI ;
  output P62ENI ;
  output P70ENI ;
  output P54ENO ;
  output P62ENO ;
  output P70ENO ;
  output P54PUON ;
  output P70PUON ;
  output P55DOUT ;
  output P63DOUT ;
  output P71DOUT ;
  output P55ENI ;
  output P63ENI ;
  output P71ENI ;
  output P55ENO ;
  output P63ENO ;
  output P71ENO ;
  output P55PUON ;
  output P71PUON ;
  output P55SELIN ;
  output P72DOUT ;
  output P72ENI ;
  output P72ENO ;
  output P72PUON ;
  output P73DOUT ;
  output P73ENI ;
  output P73ENO ;
  output P73PUON ;
  output IDADR24 ;
  output IDADR16 ;
  output P74DOUT ;
  output P74ENI ;
  output P74ENO ;
  output P74PUON ;
  output ICEDO20 ;
  output ICEDO12 ;
  output P75DOUT ;
  output P75ENI ;
  output P75ENO ;
  output P75PUON ;
  output P76DOUT ;
  output P76ENI ;
  output P76ENO ;
  output P76PUON ;
  output P77DOUT ;
  output P77ENI ;
  output P77ENO ;
  output P77PUON ;
  output PAENB ;
  output PSTN ;
  output R0A0 ;
  output MA14 ;
  output R0A1 ;
  output MA15 ;
  output R0A2 ;
  output R0A3 ;
  output R0A4 ;
  output R0A5 ;
  output R0FLAGZ ;
  output REG125ST ;
  output REGLC ;
  output REGLV ;
  output RTCCLKEN ;
  output RTRIM0 ;
  output RTRIM1 ;
  output RTRIM2 ;
  output RTRIM3 ;
  output RTRIM4 ;
  output RTRIM5 ;
  output SELIN1 ;
  output SELTAR ;
  output SRCUTCP ;
  output STOPZ ;
  output TRMCP010 ;
  output TRMCP011 ;
  output TRMCP012 ;
  output TRMCP013 ;
  output TRMCP014 ;
  output TRMRD2 ;
  output TSTN ;
  output VBRESZCP ;
  output VPBIAS ;
  output XT2ENI ;
  output VPPTS1 ;
  output VREGMV ;
  output VREGRMV ;
  output WDWR ;
  output WTRIM0 ;
  output WTRIM1 ;
  output WTRIM2 ;
  output X1ENI ;
  output X2ENI ;
  output XT1ENI ;
  output XTSTOP ;
  output XTWKUP ;
  output reg_adtyp ;
  output A19 ;
  output A18 ;
  output A17 ;
  output A16 ;
  output SELRO1 ;
  output CLKSEL1 ;
  output EXMA3 ;
  output FLSPM ;
  output EXMA1 ;
  output EXMA0 ;
  output DCE0 ;
  output DCLKSEL1 ;
  output DRDCLKC1 ;
  output DA13 ;
  output AF17 ;
  output DA12 ;
  output AF16 ;
  output SLFLASH ;
  output SVINTACK ;
  output SOFTBRK ;
  output STAGEADR1 ;
  output STAGEADR0 ;
  output SKIPEXE ;
  output PCWAITF ;
  output CPUMASK ;
  output CPUMISAL ;
  output FLREAD ;
  output IMDR10 ;
  output FLREADB3 ;
  output FLREADB2 ;
  output FLREADB1 ;
  output FLREADB0 ;
  output FCHRAM ;
  output SLMEM ;
  output SLEXM ;
  output SLBMEM ;
  output SPDEC ;
  output SPINC ;
  output SPREL ;
  output IDPOP ;
  output MDW10 ;
  output IMDR2 ;
  output CPUWR ;
  output WDOP ;
  output DMAACK ;
  output HLTST ;
  output STPST ;
  output INTACK ;
  output OCDWAIT ;
  output SVMOD ;
  output SVMODF ;
  output DRDCLK ;
  output SLDFLASH ;
  output ICEDO31 ;
  output ICEDO23 ;
  output ICEDO15 ;
  output ICEDO30 ;
  output ICEDO22 ;
  output ICEDO14 ;
  output ICEDO29 ;
  output ICEDO28 ;
  output ICEDO27 ;
  output ICEDO19 ;
  output ICEDO26 ;
  output ICEDO18 ;
  output ICEDO25 ;
  output ICEDO17 ;
  output ICEDO24 ;
  output ICEDO16 ;
  output ICEDO21 ;
  output ICEDO13 ;
  output ICEDO11 ;
  output ICEDO10 ;
  output ICEDO9 ;
  output ICEDO8 ;
  output ICEDO7 ;
  output ICEDO6 ;
  output ICEDO5 ;
  output ICEDO4 ;
  output ICEDO3 ;
  output ICEDO2 ;
  output ICEDO1 ;
  output ICEDO0 ;
  output PA19 ;
  output PC11 ;
  output PA18 ;
  output PC10 ;
  output PA17 ;
  output PA16 ;
  output PA15 ;
  output PA14 ;
  output PA9 ;
  output PC5 ;
  output PA8 ;
  output PC4 ;
  output PA7 ;
  output PC3 ;
  output PA6 ;
  output PC2 ;
  output PC19 ;
  output PC18 ;
  output PC17 ;
  output PC15 ;
  output PC14 ;
  output PC13 ;
  output PC12 ;
  output PC9 ;
  output PC8 ;
  output PC7 ;
  output PC6 ;
  output IDADR31 ;
  output IDADR23 ;
  output IDADR15 ;
  output IDADR30 ;
  output IDADR22 ;
  output IDADR14 ;
  output IDADR29 ;
  output IDADR28 ;
  output IDADR27 ;
  output IDADR19 ;
  output IDADR26 ;
  output IDADR18 ;
  output IDADR25 ;
  output IDADR17 ;
  output IDADR21 ;
  output IDADR13 ;
  output IDADR20 ;
  output IDADR12 ;
  output IDADR11 ;
  output IDADR10 ;
  output IDADR9 ;
  output IDADR8 ;
  output IDADR7 ;
  output IDADR6 ;
  output IDADR5 ;
  output IDADR4 ;
  output IDADR3 ;
  output IDADR2 ;
  output IDADR1 ;
  output IDADR0 ;
  output MA13 ;
  output MA7 ;
  output MA6 ;
  output MA5 ;
  output MA4 ;
  output MA3 ;
  output MA2 ;
  output CER ;
  output MA1 ;
  output MA0 ;
  output MDW15 ;
  output IMDR7 ;
  output MDW14 ;
  output IMDR6 ;
  output MDW13 ;
  output IMDR5 ;
  output MDW12 ;
  output IMDR4 ;
  output MDW11 ;
  output IMDR3 ;
  output MDW5 ;
  output MDW4 ;
  output MDW3 ;
  output MDW2 ;
  output MDW1 ;
  output MDW0 ;
  output EXCH ;
  output IMDR15 ;
  output IMDR14 ;
  output IMDR13 ;
  output IMDR12 ;
  output IMDR11 ;
  output IMDR9 ;
  output IMDR8 ;
  output IMDR1 ;
  output IMDR0 ;
  output RESB ;
  output FCLKRT ;
  output CIBRESRQ ;
  output FCLK1 ;
  output TMSPMD ;
  output TMBTSEL ;
  output BTFLG ;
  output READ ;
  output RDCLKP1 ;
  output SER ;
  output WED ;
  output WWR ;
  output MRG00 ;
  output MRG01 ;
  output MRG10 ;
  output MRG11 ;
  output MRG12 ;
  output PROGI ;
  output DCER ;
  output DSER ;
  output DWWR ;
  output DWED ;
  output DMRG00 ;
  output DMRG01 ;
  output DMRG10 ;
  output DMRG11 ;
  output DMRG12 ;
  output DREAD ;
  output AF19 ;
  output AF18 ;
  output AF13 ;
  output AF12 ;
  output AF11 ;
  output AF10 ;
  output AF1 ;
  output AF0 ;
  output OCDMOD ;
  output GDRAMWR ;
  output IAWRES ;
  output SVSTOPICE ;
  output SVPERI0ICE ;
  output SVPERI1ICE ;
  output MONMD ;
  output STBRELE ;
  output FRQSEL4 ;
  output R32MSTP ;
  output REQOCD ;
  output REQFL ;
  output TSELOREG ;
  output TSELIRES ;
  output TTEMP ;
  output R15KSTPZ ;
  output SYSRESB ;
  output OPLVIMDS1 ;
  output OPLVIMDS0 ;
  output SCANCLKICE ;
  output SCANMODEICE ;
  output SCANRESZICE ;
  output SCANENICE ;
  output CKSMER ;
  output TIIDER ;
  output CSPDTFLP ;
  output RAMSIZE7ICE ;
  output RAMSIZE6ICE ;
  output RAMSIZE5ICE ;
  output RAMSIZE4ICE ;
  output RAMSIZE3ICE ;
  output RAMSIZE2ICE ;
  output RAMSIZE1ICE ;
  output RAMSIZE0ICE ;
  output FLSIZE3ICE ;
  output FLSIZE2ICE ;
  output FLSIZE1ICE ;
  output FLSIZE0ICE ;
  output DFSIZE1ICE ;
  output DFSIZE0ICE ;
  output PIO00 ;
  output PIO01 ;
  output PIO02 ;
  output PIO10 ;
  output PIO03 ;
  output PIO11 ;
  output PIO04 ;
  output PIO12 ;
  output PIO20 ;
  output PIO05 ;
  output PIO13 ;
  output PIO21 ;
  output PIO06 ;
  output PIO14 ;
  output PIO22 ;
  output PIO30 ;
  output PIO15 ;
  output PIO23 ;
  output PIO31 ;
  output PIO16 ;
  output PIO24 ;
  output PIO40 ;
  output PIO17 ;
  output PIO25 ;
  output PIO41 ;
  output PIO26 ;
  output PIO42 ;
  output PIO50 ;
  output PIO27 ;
  output PIO43 ;
  output PIO51 ;
  output PIO52 ;
  output PIO60 ;
  output PIO53 ;
  output PIO61 ;
  output PIO54 ;
  output PIO62 ;
  output PIO70 ;
  output PIO55 ;
  output PIO63 ;
  output PIO71 ;
  output PIO72 ;
  output PIO73 ;
  output PIO74 ;
  output PIO75 ;
  output PIO76 ;
  output PIO77 ;
  output PIO120 ;
  output PIO121 ;
  output PIO122 ;
  output PIO130 ;
  output PIO123 ;
  output PIO124 ;
  output PIO140 ;
  output PIO137 ;
  output PIO141 ;
  output PIO146 ;
  output PIO147 ;
  output PRESADCZ ;
  output DGEN06 ;
  output DGEN05 ;
  output DGEN04 ;
  output DGEN03 ;
  output DGEN02 ;



  wire  ADEOCB ,ADSAR0 ,P52DIN ,P60DIN ,DECCER ,ADSAR1 ,P27ENI ,P43ENI ;
  wire  P51ENI ,BBMODE ,ADSAR2 ,ADSAR3 ,ADSAR4 ,ADSAR5 ,ADSAR6 ,ADSAR7 ;
  wire  P27ENO ,P43ENO ,P51ENO ,ADSAR8 ,P53DIN ,P61DIN ,ADSAR9 ,P52ENI ;
  wire  P60ENI ,DRO00 ,DRO01 ,DRO010 ,DRO011 ,DRO02 ,DRO03 ,DRO04 ;
  wire  FIHFL ,DRO05 ,DMARQ ,DRO06 ,DRO07 ,DRO08 ,GDINT ,DRO09 ;
  wire  EIRAMO0 ,EIRAMO1 ,FIHOCD ,BTBLS0 ,HVIN ,LVIOUTZNF ,MDRRAM0 ,MDRINT6 ;
  wire  MDRRAM1 ,MDRINT7 ,INTAS4C ,MDRRAM10 ,MDRRAM11 ,MDRRAM12 ,MDRRAM13 ,MDRRAM14 ;
  wire  MDRRAM15 ,MDRRAM2 ,MDRINT8 ,MDRRAM3 ,MDRINT9 ,INTAS4E ,MDRRAM4 ,MDRRAM5 ;
  wire  MDRRAM6 ,FRQSEL0 ,MDRRAM7 ,FRQSEL1 ,MDRRAM8 ,FRQSEL2 ,INTDMA0 ,MDRRAM9 ;
  wire  FRQSEL3 ,INTDMA1 ,PCLKADC ,MODE0 ,FSWE4 ,MODE1 ,FSWE5 ,OSCOUTM ;
  wire  TNFEN01 ,PSELCPU ,OSCOUTS ,TNFEN07 ,PRDRTC1 ,P00DIN ,P01DIN ,P02DIN ;
  wire  P10DIN ,P03DIN ,P11DIN ,P04DIN ,P12DIN ,P20DIN ,BBCLKR ,P05DIN ;
  wire  P13DIN ,P21DIN ,P06DIN ,P14DIN ,P22DIN ,P30DIN ,P120DIN ,P137DIN ;
  wire  P140DIN ,P141DIN ,P146DIN ,P147DIN ,P147SELIN1B5V ,P15DIN ,P23DIN ,P31DIN ;
  wire  P16DIN ,P24DIN ,P40DIN ,P17DIN ,P25DIN ,P41DIN ,BBINT0 ,P26DIN ;
  wire  P42DIN ,P50DIN ,BBINT8 ,P27DIN ,P43DIN ,P51DIN ,BBFSUB ,P40SELIN1B5V ;
  wire  P54DIN ,P62DIN ,P70DIN ,DGEN00 ,P55DIN ,P63DIN ,P71DIN ,P72DIN ;
  wire  P73DIN ,P74DIN ,P75DIN ,P76DIN ,P77DIN ,POCREL ,RESETB ,POCREL5V ;
  wire  POCRELNF ,PRDIIC14 ,R15KOUT ,R32MOUT ,RESETINBNF ,RO00 ,PID0 ,MDW6 ;
  wire  RO01 ,PID1 ,MDW7 ,MEOC ,RO010 ,PID10 ,RO011 ,PID11 ;
  wire  RO012 ,RO020 ,PID20 ,PID12 ,CPURD ,RO013 ,RO021 ,PID21 ;
  wire  PID13 ,RO014 ,RO022 ,RO030 ,PID30 ,PID22 ,PID14 ,RO110 ;
  wire  RO015 ,RO023 ,RO031 ,PID31 ,PID23 ,PID15 ,RO111 ,RO016 ;
  wire  RO024 ,RO032 ,PID24 ,PID16 ,RO120 ,RO112 ,RO017 ,RO025 ;
  wire  RO033 ,PID25 ,PID17 ,RO121 ,RO113 ,RO018 ,RO026 ,RO034 ;
  wire  PID26 ,PID18 ,RO130 ,RO122 ,RO114 ,RO019 ,RO027 ,RO035 ;
  wire  PID27 ,PID19 ,RO131 ,RO123 ,RO115 ,RO02 ,PID2 ,RO10 ;
  wire  MDW8 ,RO028 ,RO036 ,PID28 ,RO132 ,RO124 ,RO116 ,RO029 ;
  wire  RO037 ,PID29 ,RO133 ,RO125 ,RO117 ,RO03 ,PID3 ,RO11 ;
  wire  MDW9 ,RO04 ,PID4 ,RO12 ,RO05 ,PID5 ,RO13 ,RO06 ;
  wire  PID6 ,RO14 ,RO07 ,PID7 ,RO15 ,RO08 ,PID8 ,RO16 ;
  wire  EXER ,RO09 ,PID9 ,RO17 ,RPERR ,RTCCLK ,STN ,TRESET ;
  wire  VREG ,X1DIN ,RO136 ,RO128 ,EXMA2 ,X2DIN ,PER00 ,XT1DIN ;
  wire  XT2DIN ,A10 ,A11 ,A12 ,A13 ,A14 ,A15 ,A2 ;
  wire  A3 ,A4 ,A5 ,A6 ,A7 ,A8 ,A9 ,ADBIONB ;
  wire  CK0IIC0 ,ADCHSEL0 ,ADCHSEL1 ,ADCHSEL2 ,ADCHSEL3 ,ADCHSEL4 ,ADCLK ,BBMA9 ;
  wire  ADCMP ,BBFIL ,ADCPON ,ADGSELMOD ,ADINL5V ,BBHIOON ,ADOFC ,ADPDB ;
  wire  ADS1 ,ADTESMOD0 ,ADTESMOD1 ,ADTESMOD2 ,ADVSELMOD0 ,ADVSELMOD1 ,AMPH ,PC16 ;
  wire  AMPHS0 ,AMPHS1 ,AMPSEL ,BEU0 ,MA10 ,BEU1 ,MA11 ,BEU2 ;
  wire  MA12 ,BFA ,BG1ST ,BBMA0 ,BG2ADEN ,BG2ADSEL ,BGRT0 ,DFLEN ;
  wire  BGRT1 ,BGRT10 ,BGRT2 ,BGRT3 ,BGRT4 ,BGRT5 ,BGRT6 ,BGRT7 ;
  wire  BGRT8 ,BGRT9 ,BRSAM ,MDR11 ,CPUCLKEN ,CTRIM0 ,CTRIM1 ,CTRIM2 ;
  wire  CTRIM3 ,CTRIM4 ,CTRIM5 ,CTRIM6 ,DA0 ,AF2 ,DA1 ,AF3 ;
  wire  DA10 ,AF14 ,DA11 ,AF15 ,DA2 ,AF4 ,DA3 ,AF5 ;
  wire  DA4 ,CE0 ,AF6 ,DA5 ,CE1 ,AF7 ,DA6 ,AF8 ;
  wire  DA7 ,AF9 ,DA8 ,DA9 ,DSRCUT ,DTRMCP010 ,DTRMCP011 ,DTRMCP012 ;
  wire  DTRMCP013 ,DTRMCP014 ,DW0 ,MA8 ,DW1 ,MA9 ,DW10 ,DW11 ;
  wire  DW12 ,DW20 ,DW13 ,DW21 ,ALT1 ,DW14 ,DW22 ,DW30 ;
  wire  ALT2 ,DW15 ,DW23 ,DW31 ,DW16 ,DW24 ,DW32 ,DW17 ;
  wire  DW25 ,DW33 ,DDIS ,DW18 ,DW26 ,DW34 ,PA10 ,DW19 ;
  wire  DW27 ,DW35 ,PA11 ,DW2 ,DW28 ,DW36 ,PA12 ,DW29 ;
  wire  DW37 ,PA13 ,DW3 ,DW4 ,DW5 ,DW6 ,PA2 ,DW7 ;
  wire  PA3 ,DIS ,DW8 ,PA4 ,PC0 ,DW9 ,PA5 ,PC1 ;
  wire  EXA ,TA3 ,EXCLK ,EXCLKS ,FCLK2 ,FRSEL0 ,FRSEL1 ,FRSEL2 ;
  wire  FLSTOP ,FRSEL3 ,FRSEL4 ,FTRIM0 ,FTRIM1 ,FTRIM2 ,FTRIM3 ,FTRIM4 ;
  wire  FTRIM5 ,HVPPTS1 ,INCDECWS0 ,INCDECWS1 ,LOSCTEST ,LVIEN ,LVIS2 ,LVIS0 ;
  wire  LVIS1 ,LVIS3 ,LVITEST ,PSELMD2 ,LVITSEL ,TNFEN02 ,MDLYCUT ,MODENOP ;
  wire  MODERD ,MODEWR ,MSTOP ,MUTEST ,OREGSTP ,PRDMAW2 ,OSCSEL ,PREFIX ;
  wire  OSCSELS ,P00DOUT ,P00ENI ,P00ENO ,BBFCLK ,P00PUON ,BBINT2L ,P01DOUT ;
  wire  P01ENI ,P01ENO ,P01PUON ,BBINT7R ,P01SELIN ,P02DOUT ,P10DOUT ,P02ENI ;
  wire  P10ENI ,P02ENO ,P10ENO ,P02PUON ,P10PUON ,P03DOUT ,P11DOUT ,P03ENI ;
  wire  P11ENI ,P03ENO ,P11ENO ,P03PUON ,P11PUON ,P03SELIN ,P11SELIN ,P04DOUT ;
  wire  P12DOUT ,P20DOUT ,P04ENI ,P12ENI ,P20ENI ,P04ENO ,P12ENO ,P20ENO ;
  wire  P04PUON ,P12PUON ,P04SELIN ,P05DOUT ,P13DOUT ,P21DOUT ,P05ENI ,P13ENI ;
  wire  P21ENI ,P05ENO ,P13ENO ,P21ENO ,P05PUON ,P13PUON ,P06DOUT ,P14DOUT ;
  wire  P22DOUT ,P30DOUT ,P06ENI ,P14ENI ,P22ENI ,P30ENI ,P06ENO ,P14ENO ;
  wire  P22ENO ,P30ENO ,P06PUON ,P14PUON ,P30PUON ,P10SELIN ,P120DOUT ,P120ENI ;
  wire  P120ENO ,P120PUON ,P130DOUT ,P130ENO ,P137ENI ,P13SELIN ,P140DOUT ,P140ENI ;
  wire  P140ENO ,P140PUON ,P141DOUT ,P141ENI ,P141ENO ,P141PUON ,P146DOUT ,P146ENI ;
  wire  P146ENO ,P146PUON ,P147DOUT ,P147ENI ,P147ENO ,P147PUON ,P14SELIN ,P15DOUT ;
  wire  P23DOUT ,P31DOUT ,BBINT7L ,BBINT4R ,P15ENI ,P23ENI ,P31ENI ,P15ENO ;
  wire  P23ENO ,P31ENO ,P15PUON ,P31PUON ,P15SELIN ,BBREGCTL ,P16DOUT ,P24DOUT ;
  wire  P40DOUT ,P16ENI ,P24ENI ,P40ENI ,BBINT1 ,P16ENO ,P24ENO ,P40ENO ;
  wire  BBINT7 ,P16PUON ,P40PUON ,P16SELIN ,P17DOUT ,P25DOUT ,P41DOUT ,P17ENI ;
  wire  P25ENI ,P41ENI ,BBINT9 ,P17ENO ,P25ENO ,P41ENO ,P17PUON ,P41PUON ;
  wire  P17SELIN ,P26DOUT ,P42DOUT ,P50DOUT ,P26ENI ,P42ENI ,P50ENI ,P26ENO ;
  wire  P42ENO ,P50ENO ,P27DOUT ,P43DOUT ,P51DOUT ,P42PUON ,P50PUON ,P43PUON ;
  wire  P51PUON ,P52DOUT ,P60DOUT ,P52ENO ,P60ENO ,P52PUON ,P53DOUT ,P61DOUT ;
  wire  P53ENI ,P61ENI ,DGEN01 ,P53ENO ,P61ENO ,DGEN07 ,P53PUON ,P54DOUT ;
  wire  P62DOUT ,P70DOUT ,P54ENI ,P62ENI ,P70ENI ,P54ENO ,P62ENO ,P70ENO ;
  wire  P54PUON ,P70PUON ,P55DOUT ,P63DOUT ,P71DOUT ,P55ENI ,P63ENI ,P71ENI ;
  wire  P55ENO ,P63ENO ,P71ENO ,P55PUON ,P71PUON ,DMAMA12 ,P55SELIN ,P72DOUT ;
  wire  P72ENI ,P72ENO ,P72PUON ,P73DOUT ,BBRPERR ,P73ENI ,P73ENO ,P73PUON ;
  wire  IDADR24 ,IDADR16 ,P74DOUT ,P74ENI ,P74ENO ,P74PUON ,ICEDO20 ,ICEDO12 ;
  wire  P75DOUT ,P75ENI ,P75ENO ,P75PUON ,P76DOUT ,P76ENI ,P76ENO ,P76PUON ;
  wire  P77DOUT ,P77ENI ,P77ENO ,P77PUON ,PAENB ,PSTN ,R0A0 ,MA14 ;
  wire  R0A1 ,MA15 ,R0A2 ,R0A3 ,R0A4 ,R1A0 ,R0A5 ,R1A1 ;
  wire  R0FLAGZ ,REG125ST ,REGLC ,REGLV ,TIN02 ,RTCCLKEN ,RTRIM0 ,TOUT06 ;
  wire  RTRIM1 ,TOUT07 ,RTRIM2 ,RTRIM3 ,RTRIM4 ,RTRIM5 ,SELIN1 ,PRDAD5 ;
  wire  RDMRGC ,SELTAR ,SRCUTCP ,TRMCP06 ,STOPZ ,TXOCD ,TRMCP010 ,TRMCP011 ;
  wire  TRMCP012 ,TRMCP013 ,TRMCP014 ,TRMCP110 ,TRMRD2 ,TSTN ,VBRESZCP ,VPBIAS ;
  wire  XT2ENI ,VPPTS1 ,VREGMV ,VREGRMV ,WDWR ,WTRIM0 ,WTRIM1 ,WTRIM2 ;
  wire  X1ENI ,PER01 ,X2ENI ,XT1ENI ,XTSTOP ,XTWKUP ,reg_adtyp ,A19 ;
  wire  A18 ,A17 ,A16 ,SELRO1 ,CLKSEL1 ,ICETMSPMD ,ICETMBTSEL ,RO137 ;
  wire  RO129 ,EXMA3 ,FLSPM ,RO135 ,RO127 ,RO119 ,EXMA1 ,RO134 ;
  wire  RO126 ,RO118 ,EXMA0 ,RO19 ,RO18 ,DCE0 ,DCLKSEL1 ,DRDCLKC1 ;
  wire  DA13 ,AF17 ,DA12 ,AF16 ,SLFLASH ,WAITFL2 ,PRDSCN2 ,SVI ;
  wire  SVVCOUT7 ,SVVCOUT6 ,SVVCOUT5 ,SVVCOUT4 ,SVVCOUT3 ,SVVCOUT2 ,SVVCOUT1 ,SVVCOUT0 ;
  wire  SVINTACK ,SOFTBRK ,ICEMSKNMI ,ICEMSKDBG ,STAGEADR1 ,STAGEADR0 ,SKIPEXE ,PCWAITF ;
  wire  CPUMASK ,CPUPID1 ,CPUMISAL ,FLREAD ,IMDR10 ,FHLTST ,FLREADB3 ,FLREADB2 ;
  wire  FLREADB1 ,FLREADB0 ,FCHRAM ,DMAMA9 ,SLMEM ,SLEXM ,SLBMEM ,SPDEC ;
  wire  SPINC ,SPREL ,IDPOP ,MDW10 ,IMDR2 ,FLRO8 ,CPUWR ,PER04 ;
  wire  WDOP ,ICEWAITMEM ,DMAACK ,HLTST ,TID10 ,FSWS0 ,STPST ,INTACK ;
  wire  OCDWAIT ,MDRIM86 ,SVMOD ,SVMODF ,DRDCLK ,SLDFLASH ,ICECSGREGU ,ICEIFA4 ;
  wire  ICEIFA3 ,ICEIFA2 ,ICEDO31 ,ICEDO23 ,ICEDO15 ,ICEDO30 ,ICEDO22 ,ICEDO14 ;
  wire  ICEDO29 ,ICEDO28 ,ICEDO27 ,ICEDO19 ,ICEDO26 ,ICEDO18 ,ICEDO25 ,ICEDO17 ;
  wire  ICEDO24 ,ICEDO16 ,ICEDO21 ,ICEDO13 ,ICEDO11 ,DFLRO11 ,ICEDO10 ,DFLRO10 ;
  wire  ICEDO9 ,DFLRO9 ,ICEDO8 ,DETECT ,DFLRO8 ,ICEDO7 ,DFLRO7 ,ICEDO6 ;
  wire  DFLRO6 ,ICEDO5 ,DFLRO5 ,ICEDO4 ,DFLRO4 ,ICEDO3 ,DFLRO3 ,ICEDO2 ;
  wire  DFLRO2 ,ICEDO1 ,BITEN7 ,DFLRO1 ,ICEDO0 ,BITEN6 ,DFLRO0 ,PA19 ;
  wire  PC11 ,PA18 ,PC10 ,CEPR ,PA17 ,PA16 ,PA15 ,PA14 ;
  wire  PA9 ,PC5 ,PA8 ,PC4 ,PA7 ,PC3 ,PA6 ,PC2 ;
  wire  PC19 ,PC18 ,PC17 ,PC15 ,PC14 ,PC13 ,PC12 ,PC9 ;
  wire  PC8 ,PC7 ,PC6 ,IDADR31 ,IDADR23 ,IDADR15 ,IDADR30 ,IDADR22 ;
  wire  IDADR14 ,IDADR29 ,IDADR28 ,IDADR27 ,IDADR19 ,IDADR26 ,IDADR18 ,IDADR25 ;
  wire  IDADR17 ,IDADR21 ,IDADR13 ,IDADR20 ,IDADR12 ,IDADR11 ,IDADR10 ,IDADR9 ;
  wire  BITEN5 ,IDADR8 ,BITEN4 ,IDADR7 ,BITEN3 ,IDADR6 ,BITEN2 ,IDADR5 ;
  wire  BITEN1 ,IDADR4 ,BITEN0 ,IDADR3 ,IDADR2 ,IDADR1 ,IDADR0 ,MA13 ;
  wire  MA7 ,MA6 ,MA5 ,MA4 ,MA3 ,MA2 ,CER ,MA1 ;
  wire  MA0 ,MDW15 ,IMDR7 ,MDW14 ,IMDR6 ,MDW13 ,IMDR5 ,MDW12 ;
  wire  IMDR4 ,MDW11 ,IMDR3 ,FLRO9 ,MDW5 ,MDW4 ,MDW3 ,MDW2 ;
  wire  MDW1 ,MDW0 ,EXCH ,IMDR15 ,IMDR14 ,IMDR13 ,IMDR12 ,IMDR11 ;
  wire  IMDR9 ,IMDR8 ,IMDR1 ,FLRO7 ,IMDR0 ,FLRO6 ,CPUPID31 ,CPUPID23 ;
  wire  CPUPID15 ,CPUPID30 ,CPUPID22 ,CPUPID14 ,CPUPID29 ,CPUPID28 ,CPUPID27 ,CPUPID19 ;
  wire  CPUPID26 ,CPUPID18 ,CPUPID25 ,CPUPID17 ,CPUPID24 ,CPUPID16 ,CPUPID21 ,CPUPID13 ;
  wire  CPUPID20 ,CPUPID12 ,CPUPID11 ,CPUPID10 ,CPUPID9 ,CPUPID8 ,CPUPID7 ,CPUPID6 ;
  wire  FRQ4ENR ,CPUPID5 ,CPUPID4 ,CPUPID3 ,CPUPID2 ,CPUPID0 ,FRQ4ENL ,FLSIZE3 ;
  wire  FLSIZE2 ,FLSIZE1 ,FLSIZE0 ,RAMSIZE7 ,RAMSIZE6 ,RAMSIZE5 ,RAMSIZE4 ,RAMSIZE3 ;
  wire  RAMSIZE2 ,RAMSIZE1 ,RAMSIZE0 ,BFSIZE3 ,BFSIZE2 ,BFSIZE1 ,BFSIZE0 ,BMSIZE3 ;
  wire  BMSIZE2 ,BMSIZE1 ,BMSIZE0 ,DFSIZE1 ,DFSIZE0 ,ICEMKLVI ,ICEMKWDT ,ICEMKSRQ ;
  wire  RESB ,FCLKRT ,CIBRESRQ ,CIBRESRQICE ,FCLK1 ,TMSPMD ,TMBTSEL ,PRSCLK4 ;
  wire  OPWDWS0 ,BTFLG ,READ ,SP10 ,RDCLKP1 ,SER ,WED ,WWR ;
  wire  MRG00 ,MRG01 ,MRG10 ,FSWE0 ,MRG11 ,PCLK1 ,FSWE1 ,MRG12 ;
  wire  FSWE2 ,PROGI ,ICEFLERR ,ICENOECC ,DCER ,R0A6 ,R1A2 ,DSER ;
  wire  TE04 ,DWWR ,TID0 ,DWED ,TE06 ,DMRG00 ,DMRG01 ,DMRG10 ;
  wire  DMRG11 ,DMRG12 ,DREAD ,CKSEL ,AF19 ,AF18 ,AF13 ,AF12 ;
  wire  AF11 ,AF10 ,AF1 ,AF0 ,OCDMOD ,ICECK60M ,CLK60MHZ ,CLK60M ;
  wire  GDRAMWR ,IAWRES ,SVSTOPIAW ,CPUWRIAW ,PSEUDOON10 ,PSEUDOON1 ,SVSTOPICE ,SVSTOP ;
  wire  SVPERI0ICE ,SVPERI0 ,SVPERI1ICE ,SVPERI1 ,MONMD ,TOE02 ,PIOR6 ,MONSVMOD ;
  wire  STBRELE ,SOUT001 ,STBRELEICE ,FRQSEL4 ,R32MSTP ,REQOCD ,REQFL ,TSELOREG ;
  wire  TSELIRES ,TTEMP ,R15KSTPZ ,SYSRESB ,OPLVIMDS1 ,OPLVIMDS0 ,SCANCLKICE ,SCANMODEICE ;
  wire  SCANRESZICE ,SCANENICE ,SCANCLK ,SCANMODE ,SCANRESZ ,SCANEN ,FPWWR0 ,CKSMER ;
  wire  ICEDATAFLT ,ICEDMAFLT ,ICEFETCHFLT ,ICESVSTOP ,TIIDER ,PSEUDOTIIDER ,ICECKSMER ,CSPDTFLP ;
  wire  CSPDTFLG ,RAMSIZE7ICE ,RAMSIZE6ICE ,RAMSIZE5ICE ,RAMSIZE4ICE ,RAMSIZE3ICE ,RAMSIZE2ICE ,RAMSIZE1ICE ;
  wire  RAMSIZE0ICE ,FLSIZE3ICE ,FLSIZE2ICE ,FLSIZE1ICE ,FLSIZE0ICE ,DFSIZE1ICE ,DFSIZE0ICE ,SYSRSOUTB ;
  wire  PIO00 ,PCLK6 ,FSWE6 ,IREFT ,PIO01 ,FSWE7 ,PIO02 ,PIO10 ;
  wire  INTAD ,SDAI0 ,FSWE8 ,PIO03 ,PIO11 ,FSWE9 ,PIO04 ,PIO12 ;
  wire  PIO20 ,PIO05 ,PIO13 ,PIO21 ,PIO06 ,PIO14 ,PIO22 ,PIO30 ;
  wire  PIO15 ,PIO23 ,PIO31 ,PIO16 ,PIO24 ,PIO40 ,PIO17 ,PIO25 ;
  wire  PIO41 ,PIO26 ,PIO42 ,PIO50 ,PIO27 ,PIO43 ,PIO51 ,PIO52 ;
  wire  PIO60 ,INTP0 ,PIO53 ,PIO61 ,INTP1 ,PIO54 ,PIO62 ,PIO70 ;
  wire  INTP2 ,FMXST ,SDAO0 ,PIO55 ,PIO63 ,PIO71 ,INTP3 ,SDAO1 ;
  wire  PIO72 ,INTP4 ,PIO73 ,INTP5 ,PIO74 ,INTP6 ,PIO75 ,INTP7 ;
  wire  PIO76 ,INTFL ,INTP8 ,PIO77 ,INTP9 ,PIO120 ,PIO121 ,PIO122 ;
  wire  PIO130 ,PIO123 ,PIO124 ,PIO140 ,PIO137 ,PIO141 ,PIO146 ,PIO147 ;
  wire  PRESADCZ ,TESENO0L ,DGEN06 ,DGEN05 ,DGEN04 ,DGEN03 ,DGEN02 ,BBWAIT56 ;
  wire  BBWAITMEM ,MONACTIVE ,INTLVI ,INTSAU10 ,INTSAU02 ,INTSAU11 ,INTSAU03 ,INTSRE2 ;
  wire  INTSAU00 ,INTSAU01 ,INTIIC0 ,MDRPOG8 ,INTTM00 ,INTTM01 ,INTTM02 ,INTTM03 ;
  wire  INTRTC ,INTRTCI ,INTKR ,BBINT2 ,INTTM04 ,INTTM05 ,INTTM06 ,INTTM07 ;
  wire  PCLKRTC ,BBINT10 ,BBINT11 ,BBINT12 ,INTMD ,TID30 ,TID22 ,TID14 ;
  wire  FSWS4 ,BBINT13 ,BASECK ,INTSRO ,P11EXINA ,P03EXINA ,PSELCSC1 ,PSELCSC2 ;
  wire  OSCNOSTP ,TESENI2T ,PSELCSC3 ,PCLKTAU0 ,PCLKSAU0 ,MODEFNOP ,PCLKSAU1 ,PCLKIIC ;
  wire  PRESTAU0Z ,PRESSAU0Z ,PRESSAU1Z ,PRESIICZ ,PSELPOG2 ,PRESRTCZ ,PSELWWDT ,REQPCLKSAU0 ;
  wire  REQPCLKAD ,PCLKFCB ,PSELFCB1 ,PSELFCB2 ,PRDSCN10 ,PEXA ,TID9 ,SPRGMOD ;
  wire  PSELCIBC ,PSELCIB4 ,PRDSCN12 ,TESTMOD ,PRSCLK8 ,PSELCIBD ,PSELPCL ,PSELRTC ;
  wire  OPTBCT ,PRESWDTZ ,PSELMAW ,PRDRTC7 ,BASECKHS ,PSELMOD1 ,PSELMOD2 ,TR32MOUT ;
  wire  TR15KOUT ,TFIHFL ,TFIHOCD ,PRDCRC0 ,OSCOUTCP ,PRDRTC10 ,PSELOCD2 ,TIN00 ;
  wire  OTI00 ,TLVIF ,P13EXINA ,P05EXINA ,DLY50NO ,P14EXINA ,P30EXINA ,P06EXINA ;
  wire  DLY300NO ,PSELSCN ,VPPTS1_CP ,PSELPOG1 ,PSELIM8 ,P141EXINA ,P140EXINA ,INTP5EG ;
  wire  MDRMUL1 ,P31EXINA ,P15EXINA ,P51EXINA ,P43EXINA ,P50EXINA ,P42EXINA ,INTP0EG ;
  wire  PSELIM4 ,INTP11 ,INTP10 ,INTP11EG ,INTP10EG ,P75EXINA ,P74EXINA ,PSELIIC1 ;
  wire  PSELIIC2 ,SCLI0 ,SCLI1DLY ,SDAI1DLY ,PRSI000 ,PSELSA01 ,PSELSA02 ,TESENO0R ;
  wire  SEINT0SAU0 ,INTSRE0 ,SEINT2SAU0 ,INTSRE1 ,SIN03 ,SIN02 ,SIN10 ,SIN00 ;
  wire  P04EXINA ,P12EXINA ,SCKI00 ,SEL38P ,SOUT000 ,SOUT002 ,SOUT010 ,SOUT003 ;
  wire  SOUT011 ,SOUT012 ,SOUT100 ,SOUT013 ,SOUT101 ,SCKO00 ,SCKO01 ,SCKO02 ;
  wire  SCKO10 ,SCKO03 ,SCKO11 ,PCLKRW ,CK0SAU0 ,CK1SAU0 ,SNFEN00 ,PRDMAW6 ;
  wire  SNFEN10 ,TESDBT2 ,PRDMAW8 ,PRSS000 ,PRSS001 ,PRSS002 ,PRSS010 ,PRSS003 ;
  wire  PRSS011 ,PRSS012 ,PRSS100 ,PRSS013 ,PRSS101 ,PSELSA11 ,PSELSA12 ,LOWPOWER ;
  wire  TESENO1R ,TESENO0T ,SEINT0SAU1 ,P71EXINA ,P55EXINA ,P63EXINA ,P70EXINA ,P54EXINA ;
  wire  P62EXINA ,PRSS103 ,PRSS111 ,PRSS102 ,PRSS110 ,PRSS113 ,PRST001 ,PRSS112 ;
  wire  PRST000 ,SOUT110 ,SOUT111 ,CK0SAU1 ,CK1SAU1 ,SNFEN20 ,PRDPCL0 ,PSELTA01 ;
  wire  PSELTA02 ,INTTM01H ,INTTM03H ,CKENTAU07 ,CKENTAU06 ,CKENTAU05 ,CKENTAU04 ,CKENTAU03 ;
  wire  CKENTAU02 ,CKENTAU01 ,CKENTAU00 ,TOUT00 ,TOUT01 ,TOUT02 ,TOUT03 ,TOUT04 ;
  wire  TOUT05 ,TIN07O ,MONPC7 ,PRDAD1 ,TIN06 ,TIN05O ,MONPC3 ,TIN04 ;
  wire  TDIN4 ,TIN03 ,TDIN3 ,P16EXINA ,TE07 ,TE05 ,TE03 ,TE02 ;
  wire  TE01 ,TE00 ,TOE07 ,TOE06 ,TOE05 ,TOE04 ,TOE03 ,PIOR7 ;
  wire  TOE01 ,PIOR5 ,TOE00 ,PIOR4 ,PRST002 ,PRST010 ,PRST003 ,PRST011 ;
  wire  PRST012 ,PRST020 ,OPWDINT ,PRST013 ,PRST021 ,PRST030 ,PRST031 ,TNFEN00 ;
  wire  TNFEN03 ,TNFEN04 ,TNFEN05 ,TNFEN06 ,PRDRTC0 ,CK0TAU0 ,CK1TAU0 ,CK2TAU0 ;
  wire  BBINT1L ,CK3TAU0 ,BBINT9L ,BBINT6R ,SOUT012DLY ,SOUT010DLY ,SOUT011DLY ,SOUT013DLY ;
  wire  SOUT110DLY ,SOUT111DLY ,PSELAD1 ,PRDMAW3 ,PSELAD2 ,PRDMAW4 ,ADTRIG0 ,PSELP0 ;
  wire  PRDP0000 ,PRDP0001 ,PRDP0002 ,PRDP0003 ,PRDP0004 ,PRDP0005 ,PRDP0006 ,PRDP0110 ;
  wire  PRDP0007 ,PRDP0111 ,P00EXOUTA ,P00EXINA ,P01EXOUTB ,P01EXINA ,P02EXOUTA ,P10EXOUTA ;
  wire  P02EXINA ,P10EXINA ,P03EXOUTB ,P11EXOUTB ,P05EXOUTB ,P13EXOUTB ,P06EXOUTB ,P14EXOUTB ;
  wire  PORT0EXOR ,PSELP1 ,PRDP0108 ,PRDP0204 ,PRDP0109 ,PRDP0205 ,PRDP0112 ,PRDP0200 ;
  wire  PRDP0113 ,PRDP0201 ,PRDP0114 ,PRDP0202 ,PRDP0115 ,PRDP0203 ,P10EXOUTB ,P10EXOUTC ;
  wire  P11EXOUTC ,P12EXOUTB ,P13EXOUTA ,P13EXOUTC ,P14EXOUTC ,P15EXOUTB ,P31EXOUTB ,P15EXOUTC ;
  wire  P31EXOUTC ,P16EXOUTA ,P17EXOUTA ,P17EXOUTB ,P41EXOUTB ,P17EXINA ,P41EXINA ,PORT1EXOR ;
  wire  P10EXINB ,P12EXINB ,BBINT11L ,PSELP2 ,PRES6Z ,PRDP0206 ,PRDP0310 ,MONMDW10 ;
  wire  PRDP0207 ,PRDP0311 ,MONMDW11 ,PORT2EXOR ,PSELP3 ,PRDP0308 ,PRDP0404 ,PRDP1204 ;
  wire  PRDP0309 ,PRDP0405 ,PRDP1205 ,PRDP0312 ,PRDP0400 ,PRDP1200 ,MONMDW12 ,PRDP0313 ;
  wire  PRDP0401 ,PRDP1201 ,MONMDW13 ,PRDP0314 ,PRDP0402 ,PRDP1202 ,MONMDW14 ,PRDP0315 ;
  wire  PRDP0403 ,PRDP1203 ,MONMDW15 ,CLK1HZ ,PORT3EXOR ,PSELP4 ,PRDP0406 ,PRDP0510 ;
  wire  PRDP1206 ,PRDP1310 ,PRDP0407 ,PRDP0511 ,PRDP1207 ,PRDP1311 ,P42EXOUTB ,PORT4EXOR ;
  wire  PSELP5 ,PRDP0508 ,PRDP0604 ,PRDP1308 ,PRDP1404 ,PRDP0509 ,PRDP0605 ,PRDP1309 ;
  wire  PRDP1405 ,PRDP0512 ,PRDP0600 ,PRDP1312 ,PRDP1400 ,PRDP0513 ,PRDP0601 ,PRDP1313 ;
  wire  PRDP1401 ,PRDP0514 ,PRDP0602 ,PRDP1314 ,PRDP1402 ,PRDP0515 ,PRDP0603 ,PRDP1315 ;
  wire  PRDP1403 ,P51EXOUTA ,P52EXINA ,P60EXINA ,P53EXINA ,P61EXINA ,P55EXOUTA ,P55EXOUTB ;
  wire  PORT5EXOR ,PSELP6 ,PRDP0606 ,PRDP0710 ,PRDP1406 ,PRDP0607 ,PRDP0711 ,PRDP1407 ;
  wire  P60EXOUTB ,P61EXOUTB ,PORT6EXOR ,PSELP7 ,PRDP0708 ,PRDP0709 ,PRDP0712 ,PRDP0713 ;
  wire  PRDP0714 ,PRDP0715 ,P72EXINA ,P73EXINA ,P76EXINA ,BBPWRITE ,P77EXOUTA ,P77EXINA ;
  wire  PORT7EXOR ,PSELP12 ,PRDMOD8 ,P120EXINA ,P122EXINA ,PORT12EXOR ,PSELP13 ,PRDMOD9 ;
  wire  P137EXINA ,PSELP14 ,P140EXOUTB ,P141EXOUTB ,P146EXINA ,P147EXINA ,PORT14EXOR ,BBREQPCLKL ;
  wire  BBCKSELRL ,BBCKSELML ,BBHIOONL ,BBREGCTLL ,BBPRDATA15L ,BBPRDATA12R ,BBPRDATA14L ,BBPRDATA11R ;
  wire  BBPRDATA13L ,BBPRDATA10R ,BBPRDATA12L ,BBPRDATA11L ,BBPRDATA10L ,BBPRDATA9L ,BBPRDATA6R ,BBPRDATA8L ;
  wire  BBPRDATA5R ,BBPRDATA7L ,BBPRDATA4R ,BBPRDATA6L ,BBPRDATA3R ,BBPRDATA5L ,BBPRDATA2R ,BBPRDATA4L ;
  wire  BBPRDATA1R ,BBPRDATA3L ,BBPRDATA0R ,BBPRDATA2L ,BBPRDATA1L ,BBPRDATA0L ,BBWAITMEML ,BBWAIT56L ;
  wire  BBINT0L ,BBINT3L ,BBINT0R ,BBINT4L ,BBINT1R ,BBINT5L ,BBINT2R ,BBINT6L ;
  wire  BBINT3R ,BBINT8L ,BBINT5R ,BBINT10L ,BBINT12L ,BBINT13L ,BBINT10R ,BBMODEL ;
  wire  BBSCANOUTL ,ADTRIG0L ,ADTRIG1L ,INTRTDISL ,BBCLKRL ,BBFMAIN ,BBCLKML ,TESSCAN1 ;
  wire  BBREQPCLKR ,BBCKSELRR ,BBCKSELMR ,BBHIOONR ,BBREGCTLR ,BBPRDATA15R ,BBPRDATA14R ,BBPRDATA13R ;
  wire  BBPRDATA9R ,BBPRDATA8R ,BBPRDATA7R ,BBWAITMEMR ,BBWAIT56R ,BBINT8R ,BBINT9R ,BBINT11R ;
  wire  BBINT12R ,BBINT13R ,BBMODER ,BCKHSEN ,BBSCANOUTR ,ADTRIG0R ,ADTRIG1R ,INTRTDISR ;
  wire  BBCLKRR ,BBCLKMR ,pull_down0 ,pull_down1 ,pull_down2 ,pull_down3 ,pull_down4 ,pull_down5 ;
  wire  pull_down6 ,pull_down7 ,pull_down8 ,pull_down9 ,pull_down10 ,pull_down11 ,pull_down12 ,pull_down20 ;
  wire  pull_down13 ,pull_down21 ,pull_down14 ,pull_down22 ,pull_down30 ,pull_down15 ,pull_down23 ,pull_down31 ;
  wire  pull_down16 ,pull_down24 ,pull_down32 ,pull_down40 ,pull_down17 ,pull_down25 ,pull_down33 ,pull_down41 ;
  wire  pull_down18 ,pull_down26 ,pull_down34 ,pull_down42 ,pull_down50 ,pull_down19 ,pull_down27 ,pull_down35 ;
  wire  pull_down43 ,pull_down51 ,pull_down28 ,pull_down36 ,pull_down44 ,pull_down52 ,pull_down60 ,pull_down29 ;
  wire  pull_down37 ,pull_down45 ,pull_down53 ,pull_down61 ,pull_down38 ,pull_down46 ,pull_down54 ,pull_down62 ;
  wire  pull_down70 ,pull_down39 ,pull_down47 ,pull_down55 ,pull_down63 ,pull_down71 ,pull_down48 ,pull_down56 ;
  wire  pull_down64 ,pull_down72 ,pull_down80 ,pull_down49 ,pull_down57 ,pull_down65 ,pull_down73 ,pull_down81 ;
  wire  pull_down58 ,pull_down66 ,pull_down74 ,pull_down82 ,pull_down90 ,pull_down59 ,pull_down67 ,pull_down75 ;
  wire  pull_down83 ,pull_down91 ,pull_down68 ,pull_down76 ,pull_down84 ,pull_down92 ,pull_down69 ,pull_down77 ;
  wire  pull_down85 ,pull_down93 ,pull_down78 ,pull_down86 ,pull_down94 ,pull_down79 ,pull_down87 ,pull_down95 ;
  wire  pull_down88 ,pull_down96 ,pull_down89 ,pull_down97 ,pull_down98 ,pull_down99 ,pull_down100 ,pull_down101 ;
  wire  pull_down102 ,pull_down110 ,pull_down103 ,pull_down111 ,pull_down104 ,pull_down112 ,pull_down120 ,pull_down105 ;
  wire  pull_down113 ,pull_down106 ,pull_down114 ,pull_down107 ,pull_down115 ,pull_down108 ,pull_down116 ,pull_down109 ;
  wire  pull_down117 ,pull_down118 ,pull_down119 ,pull_up0 ,pull_up1 ,pull_up2 ,pull_up3 ,pull_up4 ;
  wire  pull_up5 ,pull_up6 ,pull_up7 ,pull_up8 ,pull_up9 ,pull_up10 ,pull_up11 ,pull_up12 ;
  wire  pull_up20 ,pull_up13 ,pull_up21 ,pull_up14 ,pull_up22 ,pull_up30 ,pull_up15 ,pull_up23 ;
  wire  pull_up31 ,pull_up16 ,pull_up24 ,pull_up32 ,pull_up40 ,pull_up17 ,pull_up25 ,pull_up33 ;
  wire  pull_up41 ,pull_up18 ,pull_up26 ,pull_up34 ,pull_up42 ,pull_up50 ,pull_up19 ,pull_up27 ;
  wire  pull_up35 ,pull_up43 ,pull_up51 ,pull_up28 ,pull_up36 ,pull_up44 ,pull_up52 ,pull_up60 ;
  wire  pull_up29 ,pull_up37 ,pull_up45 ,pull_up53 ,pull_up61 ,pull_up38 ,pull_up46 ,pull_up54 ;
  wire  pull_up62 ,pull_up70 ,pull_up39 ,pull_up47 ,pull_up55 ,pull_up63 ,pull_up71 ,pull_up48 ;
  wire  pull_up56 ,pull_up64 ,pull_up72 ,pull_up49 ,pull_up57 ,pull_up65 ,pull_up73 ,pull_up58 ;
  wire  pull_up66 ,pull_up74 ,pull_up59 ,pull_up67 ,pull_up75 ,pull_up68 ,pull_up76 ,pull_up69 ;
  wire  pull_up77 ,pull_up78 ,pull_up79 ,MDRINT15 ,MDRINT14 ,MDRINT13 ,MDRINT12 ,MDRINT11 ;
  wire  MDRINT10 ,MDRINT5 ,INTAS4A ,MDRINT4 ,MDRINT3 ,MDRINT2 ,MDRINT1 ,MDRINT0 ;
  wire  MDRDMA15 ,MDRDMA14 ,MDRDMA13 ,MDRDMA12 ,MDRDMA11 ,MDRDMA10 ,MDRDMA9 ,MDRDMA8 ;
  wire  MDRDMA7 ,MDRDMA6 ,MDRDMA5 ,MDRDMA4 ,MDRDMA3 ,MDRDMA2 ,MDRDMA1 ,MDRDMA0 ;
  wire  MDRMUL15 ,MDRMUL14 ,MDRMUL13 ,MDRMUL12 ,MDRMUL11 ,MDRMUL10 ,MDRMUL9 ,PENABLE ;
  wire  MDRMUL8 ,MDRMUL7 ,MDRMUL6 ,MDRMUL5 ,PCLBUZ1 ,SEL24PI ,SEL32PI ,SEL40PI ;
  wire  MDRMUL4 ,PCLBUZ0 ,MDRMUL3 ,MDRMUL2 ,MDRMUL0 ,MDROCD15 ,MDROCD14 ,MDROCD13 ;
  wire  MDROCD12 ,MDROCD11 ,MDROCD10 ,MDROCD9 ,MDROCD8 ,MDROCD7 ,MDROCD6 ,MDROCD5 ;
  wire  MDROCD4 ,MDROCD3 ,MDROCD2 ,MDROCD1 ,MDROCD0 ,PRDCSC15 ,PRDCSC14 ,PRDCSC13 ;
  wire  PRDCSC12 ,PRDCSC11 ,PRDCSC10 ,PRDCSC9 ,PRDIIC1 ,PRDCSC8 ,PRDIIC0 ,RDSETUP ;
  wire  PRDCSC7 ,PRDCSC6 ,PRDCSC5 ,PRDCRC9 ,PRDCSC4 ,PRDCRC8 ,PRDCSC3 ,PRDCRC7 ;
  wire  PRDCSC2 ,PRDCRC6 ,PRDCSC1 ,PRDCRC5 ,PRDCSC0 ,PRDCRC4 ,PRDFCB15 ,PRDCIC11 ;
  wire  PRDFCB14 ,PRDCIC10 ,PRDFCB13 ,PRDFCB12 ,PRDFCB11 ,PRDFCB10 ,PRDFCB9 ,PRDCIC7 ;
  wire  PRDCID5 ,PRDFCB8 ,PRDCIC6 ,PRDCID4 ,PRDFCB7 ,PRDCIC5 ,PRDCID3 ,PRDFCB6 ;
  wire  PRDCIC4 ,PRDCID2 ,PRDFCB5 ,PRDCIC3 ,PRDCID1 ,PRDFCB4 ,PRDCIC2 ,PRDCID0 ;
  wire  PRDFCB3 ,PRDCIC1 ,PRDFCB2 ,PRDCIC0 ,PRDFCB1 ,RT0MON1 ,PRDFCB0 ,RT0MON0 ;
  wire  PRDCIC15 ,PRDCID11 ,PRDCIC14 ,PRDCID10 ,PRDCIC13 ,PRDCIC12 ,PRDCIC9 ,PRDCID7 ;
  wire  PRDCIC8 ,PRDCID6 ,PRDCID15 ,PRDCID14 ,PRDCID13 ,PRDCID12 ,PRDCID9 ,PRDCID8 ;
  wire  MDRCID15 ,MDRCID14 ,MDRCID13 ,MDRCID12 ,MDRCID11 ,MDRCID10 ,MDRCID9 ,MDRCID8 ;
  wire  MDRCID7 ,MDRCID6 ,MDRCID5 ,MDRCID4 ,MDRCID3 ,MDRCID2 ,MDRCID1 ,MDRCID0 ;
  wire  PRDPCL15 ,PRDPCL11 ,PRDPCL10 ,PRDPCL9 ,PRDMOD1 ,PRDPCL8 ,PRDMOD0 ,PRDPCL7 ;
  wire  PRDPCL3 ,PRDPCL2 ,PRDPCL1 ,PRDRTC15 ,PRDRTC14 ,PRDRTC13 ,PRDRTC12 ,PRDSELEN ;
  wire  OSCOUTEN ,PRDRTC11 ,PRDRTC9 ,PRDRTC8 ,PRDRTC6 ,PRDRTC5 ,WAITMEM ,PRDRTC4 ;
  wire  PRDRTC3 ,PRDRTC2 ,PRDWDT15 ,PRDWDT12 ,PRDWDT11 ,PRDWDT9 ,PRDMAW15 ,PRDMAW14 ;
  wire  PRDMAW13 ,PRDMAW12 ,PRDMAW11 ,PRDMAW10 ,PRDMAW9 ,PRDMAW7 ,PRDMAW5 ,PRDMAW1 ;
  wire  PRDMAW0 ,MONMA15 ,MONMA14 ,MONMA13 ,MONMA12 ,MONMA11 ,MONMA10 ,MONMA9 ;
  wire  RDMRG1 ,MONMA8 ,RDMRG0 ,MONMA7 ,MONMA6 ,MONMA5 ,MONMA4 ,MONMA3 ;
  wire  MONMA2 ,MONMA1 ,MONMA0 ,TDIN2B ,MONPC19 ,MONPC18 ,MONPC17 ,MONPC16 ;
  wire  MONPC15 ,MONPC14 ,MONPC13 ,MONPC12 ,MONPC11 ,MONPC10 ,MONPC9 ,PRDAD3 ;
  wire  MONPC8 ,PRDAD2 ,MONPC6 ,PRDAD0 ,MONPC5 ,MONPC4 ,MONPC2 ,TDIN2T ;
  wire  MONPC1 ,MONPC0 ,TDIN2R ,TDIN1T ,PRDCRC15 ,PRDCRC14 ,PRDCRC13 ,PRDCRC12 ;
  wire  PRDCRC11 ,PRDCRC10 ,PRDCRC3 ,PRDCRC2 ,PRDCRC1 ,PRDMOD15 ,PRDMOD14 ,PRDMOD13 ;
  wire  PRDMOD12 ,PRDMOD11 ,PRDMOD10 ,PRDMOD7 ,PRDMOD6 ,PSELBCD ,PRDMOD5 ,PRDMOD4 ;
  wire  PRDMOD3 ,PRDMOD2 ,PRDSCN15 ,PRDSCN14 ,PRDSCN13 ,PRDSCN11 ,PRDSCN9 ,PRDSCN8 ;
  wire  PRDSCN7 ,PRDSCN6 ,TESENI4 ,PRDSCN5 ,TESENI3 ,PRDSCN4 ,PRDSCN3 ,PRDSCN1 ;
  wire  PRDSCN0 ,TRMCP00 ,TSELBGR ,TRMCP01 ,TRMCP02 ,TRMCP03 ,TRMCP04 ,TRMCP05 ;
  wire  TRMCP07 ,TRMCP08 ,TRMCP09 ,TRMCP015 ,TRMCP111 ,TRMCP016 ,TRMCP112 ,TRMCP017 ;
  wire  TRMCP113 ,RTRMCP015 ,RTRMCP016 ,RTRMCP017 ,RTRMCP018 ,RTRMCP019 ,RTRMCP020 ,MDRPOG15 ;
  wire  MDRPOG14 ,MDRPOG13 ,MDRPOG12 ,MDRPOG11 ,MDRPOG10 ,MDRPOG9 ,MDRPOG7 ,SEL30PI ;
  wire  MDRPOG6 ,MDRPOG5 ,MDRPOG4 ,MDRPOG3 ,MDRPOG2 ,MDRPOG1 ,MDRPOG0 ,MDRIM815 ;
  wire  MDRIM814 ,MDRIM813 ,MDRIM812 ,MDRIM811 ,MDRIM810 ,MDRIM89 ,MDRIM88 ,MDRIM87 ;
  wire  MDRIM85 ,MDRIM84 ,MDRIM83 ,IONCHK1 ,MDRIM82 ,MDRIM81 ,MDRIM49 ,MDRIM80 ;
  wire  MDRIM48 ,MDRIM411 ,MDRIM410 ,MDRIM43 ,MDRIM42 ,MDRIM41 ,MDRIM40 ,PRDIIC15 ;
  wire  PRDIIC13 ,PRDIIC12 ,PRDIIC11 ,PRDIIC10 ,SLECCOFF ,PRDIIC9 ,PRDIIC8 ,TDSEL0B ;
  wire  PRDIIC7 ,PRDIIC6 ,PRDIIC5 ,PRDIIC4 ,PRDIIC3 ,PRDIIC2 ,PRDSA015 ,PRDSA111 ;
  wire  PRDSA014 ,PRDSA110 ,PRDSA013 ,PRDSA012 ,PRDSA011 ,PRDSA010 ,PRDSA09 ,PRDSA17 ;
  wire  PRDTA01 ,PRDSA08 ,PRDSA16 ,PRDTA00 ,TDSEL0L ,PRDSA07 ,PRDSA15 ,PRDSA06 ;
  wire  PRDSA14 ,PRDSA05 ,PRDSA13 ,PRDSA04 ,PRDSA12 ,OPOCDEN ,PRDSA03 ,PRDSA11 ;
  wire  PRDSA02 ,PRDSA10 ,TDSEL2B ,PRDSA01 ,PRDSA00 ,TDSEL1B ,PRDSA115 ,PRDSA114 ;
  wire  PRDSA113 ,PRDSA112 ,PRDSA19 ,PRDTA03 ,PRDSA18 ,PRDTA02 ,TDSEL1L ,PRDTA015 ;
  wire  PRDTA014 ,PRDTA013 ,PRDTA012 ,PRDTA011 ,PRDTA010 ,PRDTA09 ,PRDTA08 ,TDSEL1R ;
  wire  TDSEL0T ,PRDTA07 ,PRDTA06 ,TDSEL0R ,PRDTA05 ,PRDTA04 ,TDSEL2L ,PRDAD15 ;
  wire  PRDAD14 ,PRDAD13 ,PRDAD12 ,PRDAD11 ,PRDAD10 ,PRDAD9 ,PRDAD8 ,OPBOEN ;
  wire  PRDAD7 ,PRDAD6 ,PRDAD4 ,DMAMA15 ,DMAMA14 ,DMAMA13 ,DMAMA11 ,DMAMA10 ;
  wire  DMAMA8 ,DMAMA7 ,DMAMA6 ,DMAMA5 ,DMAMA4 ,DMAMA3 ,DMAMA2 ,DMAMA1 ;
  wire  DMAMA0 ,DMARD ,DMAWR ,FMAIN ,DMAWDOP ,DMAEN ,SLIRAM ,STBEN ;
  wire  MDR15 ,MDR14 ,MDR13 ,MDR12 ,IAWEN ,MDR10 ,MDR9 ,MDR8 ;
  wire  MDR7 ,MDR6 ,BTPR ,MDR5 ,MDR4 ,MDR3 ,MDR2 ,MDR1 ;
  wire  MDR0 ,VCOUT6 ,VCOUT5 ,VCOUT4 ,VCOUT3 ,OPTRAM ,VCOUT2 ,VCOUT1 ;
  wire  INTDBG ,INTNMI ,INTRQ1 ,INTRQ3 ,INTRQ2 ,INTRQ0 ,MONMDSTP ,BRKMSK ;
  wire  WAITMOD ,DMAWAIT ,SP15 ,SP14 ,FSPR ,SP13 ,SP12 ,MEOR ;
  wire  SP11 ,SP9 ,SP8 ,RDT ,SP7 ,SP6 ,SP5 ,SP4 ;
  wire  SP3 ,SP2 ,SP1 ,SP0 ,CPUSTART ,GOFIRM ,PADDR1 ,MONMDR15 ;
  wire  MONMDR14 ,MONMDR13 ,MONMDR12 ,MONMDR11 ,MONMDR10 ,MONMDR9 ,MONMDR8 ,MONMDR7 ;
  wire  MONMDR6 ,MONMDR5 ,MONMDR4 ,MONMDR3 ,MONMDR2 ,MONMDR1 ,MONMDR0 ,MONMDW9 ;
  wire  MONMDW8 ,MONMDW7 ,MONMDW6 ,MONMDW5 ,MONMDW4 ,MONMDW3 ,MONMDW2 ,MONMDW1 ;
  wire  MONMDW0 ,CRCHLTEN ,INTAS02 ,INTAS04 ,INTAS22 ,INTAS50 ,INTAS28 ,INTAS52 ;
  wire  INTAS54 ,PSELINT1 ,PSELDMAC ,PSELMD1 ,PRESOCDZ ,PCLKOCD ,OCDRESMK ,RXOCD ;
  wire  PSELOCD1 ,OCDASEN ,SLTRXTX ,OPWDEN ,GDRAM1 ,GDRAM0 ,PADDR2 ,PADDR0 ;
  wire  PWRITE ,OPTIDDQ ,OPLVIS1 ,OPLVIS0 ,EXCLK1 ,NVMRCEND ,TESSCAN3 ,TESSCAN4 ;
  wire  OPWDSTBY ,PTESINST ,TESUSR ,TESDBT ,PRES1Z ,OPTEXCCK ,WDTRES ,NSRESB ;
  wire  RESSTP ,RESSQSTA ,FSTPST ,PSUBMODE ,TPOCREL ,SRESREQ ,TFLSTOPC ,TFLSTOPD ;
  wire  PER07 ,PER06 ,PER05 ,PER03 ,PER02 ,STPBCKBT ,BBCKSELR ,BBCKSELM ;
  wire  PRSCLK1 ,VCPRGWE ,PRSCLK2 ,PRSCLK3 ,PRSCLK5 ,OPWDWS1 ,PRSCLK6 ,PRSCLK7 ;
  wire  PRSCLK9 ,PRSCLK10 ,OPTMDUMP ,PRSCLK11 ,PRSCLK12 ,PRSCLK13 ,PRSCLK14 ,PRSCLK15 ;
  wire  RT0LPM ,TMDENCLK ,BBCLKM ,INCDECMD ,BBREQPCLK ,INTRCLK ,WDTTESCK ,PCLKTST ;
  wire  SBRFONLY ,FSUB ,STDWAIT ,HISPEED ,HIOMSK ,RLOWSPY ,OPVPOC2 ,OPVPOC1 ;
  wire  OPVPOC0 ,FLROACT ,EEEMD ,WDEN ,MCM0 ,RSTS ,REQR32M ,VSETEND ;
  wire  BBCKSTR ,PSYSRESB ,BBCKSTM ,GOFIRMR ,SUBCKST ,TRMRD1 ,PADDR3 ,OPWDCS1 ;
  wire  OPWDCS0 ,PORTSELB ,OPWDCS2 ,C3HFF ,FLRO37 ,FLRO29 ,FLRO36 ,FLRO28 ;
  wire  FLRO35 ,FLRO27 ,FLRO19 ,FLRO34 ,FLRO26 ,FLRO18 ,FLRO33 ,FLRO25 ;
  wire  FLRO17 ,FLRO32 ,FLRO24 ,FLRO16 ,FLRO31 ,FLRO23 ,FLRO15 ,FLRO30 ;
  wire  FLRO22 ,FLRO14 ,FLRO21 ,FLRO13 ,FLRO20 ,FLRO12 ,FLRO11 ,FLRO10 ;
  wire  FLRO5 ,FLRO4 ,FLRO3 ,FLRO2 ,FLRO1 ,FLRO0 ,SACEEN ,EXCHEN ;
  wire  SECEN ,FSWEN ,TID20 ,TID12 ,FSWS2 ,TRMCP114 ,SRCUT ,SUB ;
  wire  TID31 ,TID23 ,TID15 ,FSWS5 ,TID29 ,TID28 ,TID27 ,TID19 ;
  wire  FSWS9 ,TID26 ,TID18 ,FSWS8 ,TID25 ,TID17 ,FSWS7 ,TID24 ;
  wire  TID16 ,FSWS6 ,TID21 ,TID13 ,FSWS3 ,TID11 ,FSWS1 ,TID8 ;
  wire  TID7 ,TID6 ,TID5 ,TID4 ,TID3 ,TID2 ,TID1 ,TESINST ;
  wire  BBTESINST ,OPTFLMEM ,TA17 ,TA16 ,TA15 ,TA14 ,TA13 ,TA12 ;
  wire  TA11 ,TA10 ,TA9 ,TA8 ,TA7 ,TA6 ,TA5 ,TA4 ;
  wire  TA2 ,TA1 ,TA0 ,TPIDSEL ,BBNVM1 ,BBNVM2 ,CFNSD9 ,CFNSD8 ;
  wire  CFNSD7 ,CFNSD6 ,CFNSD5 ,CFNSD4 ,CFNSD3 ,CFNSD2 ,CFNSD1 ,CFNSD0 ;
  wire  FSWE3 ,SELTAF ,CECCE ,TRMRD1CK ,TRMRD2CK ,RDPR ,WRPR ,SEPR ;
  wire  BTBLS1 ,FPSER2 ,FPSER1 ,FPSER0 ,FPWWR2 ,FPWWR1 ,FPERTY7 ,FPERTY6 ;
  wire  FPERTY5 ,FPERTY4 ,FPERTY3 ,FPERTY2 ,FPERTY1 ,FPERTY0 ,FPWRTY7 ,FPWRTY6 ;
  wire  FPWRTY5 ,FPWRTY4 ,FPWRTY3 ,FPWRTY2 ,FPWRTY1 ,FPWRTY0 ,FPECC3 ,FPECC2 ;
  wire  FPECC1 ,FPECC0 ,R1FLAGZ ,R0A7 ,R1A3 ,R1A7 ,R1A6 ,R1A5 ;
  wire  R1A4 ,ECCER ,FMULTIEN ,POSCNOST ,POSCOUTE ,CPT ,TESTRMRD ,AisRSEQ ;
  wire  FRQ4EN ,CHMOD ,SELTADF ,DFLSTOP ,DECCE ,OPTDFL ,LOWSPY ,CWEE ;
  wire  PADDR4 ,FLMEMTES ,MSWR ,STCHK ,WDT1 ,WDT2 ,WDT3 ,WDT4 ;
  wire  CPBT ,EXTVPP2 ,EXTVPP1 ,MODIDIS ,VCEQ ,INTWWDT ,WDTMON ,PSELCRC ;
  wire  TESSCAN2 ,OPTOPLRD ,RAMMULTI ,RAEDIS ,STAYTES ,LFSSCAIN ,TDIN5 ,TIN05 ;
  wire  TDIN1R ,TDIN0T ,TDIN1B ,TDIN0R ,TDIN0B ,TESENI2R ,TESENI1T ,TESENI2B ;
  wire  TESENI2L ,TESENI1R ,TESENI0T ,TESENI1B ,TESENI1L ,TESENI0R ,TESENI0B ,TESENI0L ;
  wire  TESENO3 ,TESENO2T ,TESENO2R ,TESENO1T ,TESENO2B ,TESENO2L ,TESENO1B ,TESENO1L ;
  wire  TESENO0B ,TDSEL3 ,TDSEL2T ,TDSEL2R ,TDSEL1T ,TDOUT3 ,TDOUT2 ,TDOUT1 ;
  wire  TDOUT0 ,SCANIN ,SCANENMD ,BBSCANOUT ,RDCLKC1 ,FLREGENB ,VCPHV ,BBPRDATA15 ;
  wire  BBPRDATA14 ,BBPRDATA13 ,BBPRDATA12 ,BBPRDATA11 ,BBPRDATA10 ,BBPRDATA9 ,BBPRDATA8 ,BBPRDATA7 ;
  wire  BBPRDATA6 ,BBPRDATA5 ,BBPRDATA4 ,BBPRDATA3 ,BBPRDATA2 ,BBPRDATA1 ,BBPRDATA0 ,BBPENABLE ;
  wire  BBMA15 ,BBMA14 ,BBMA13 ,BBMA12 ,BBMA11 ,BBMA10 ,BBMA8 ,BBMA7 ;
  wire  BBMA6 ,BBMA5 ,BBMA4 ,BBMA3 ,BBMA2 ,BBMA1 ,PADDR6 ,PADDR5 ;
  wire  PSELKR ,BBSELSFR1 ,BBSELSFR2 ,SLAPB ,MDWFLRO15 ,MDWFLRO14 ,MDWFLRO13 ,MDWFLRO12 ;
  wire  MDWFLRO11 ,MDWFLRO10 ,MDWFLRO9 ,MDWFLRO8 ,MDWFLRO7 ,MDWFLRO6 ,MDWFLRO5 ,MDWFLRO4 ;
  wire  MDWFLRO3 ,MDWFLRO2 ,MDWFLRO1 ,MDWFLRO0 ,GDPORT ,GDCSC ,TIN07 ,PIOR3 ;
  wire  PIOR2 ,PIOR1 ,PIOR0 ,SEL20P ,SEL24P ,SEL32P ,SEL40P ,SEL08P ;
  wire  SEL30P ,SEL36P ,SEL44P ,SEL52P ,SEL48P ,SEL64P ,SEL20PI ,SEL36PI ;
  wire  SEL44PI ,SEL52PI ,SEL38PI ,SEL48PI ,SEL64PI ,BBISC ,BBINT3 ,BBINT4 ;
  wire  BBINT5 ,BBINT6 ,SCLO0 ,SCLO1 ,CDEN7 ,CDEN6 ,CDEN5 ,CDEN4 ;
  wire  CDEN3 ,CDEN2 ,CDEN1 ,CDEN0 ,TXSAU ,BBSFDIS1 ,BBEXAD10 ,BBEXAD11 ;
  wire  BBEXAD12 ,BBEXOR10 ,BBEXOR11 ,BBEXOR12 ,BBSWPPT1 ,BBSWPICA ,TTRG2 ,BBMOSC ;
  wire  BBHIOSC ,ADINLBB5V ;


  TBCLL pulldown0 ( pull_down0 ) ;
  TBCLL pulldown1 ( pull_down1 ) ;
  TBCLL pulldown2 ( pull_down2 ) ;
  TBCLL pulldown3 ( pull_down3 ) ;
  TBCLL pulldown4 ( pull_down4 ) ;
  TBCLL pulldown5 ( pull_down5 ) ;
  TBCLL pulldown6 ( pull_down6 ) ;
  TBCLL pulldown7 ( pull_down7 ) ;
  TBCLL pulldown8 ( pull_down8 ) ;
  TBCLL pulldown9 ( pull_down9 ) ;
  TBCLL pulldown10 ( pull_down10 ) ;
  TBCLL pulldown11 ( pull_down11 ) ;
  TBCLL pulldown12 ( pull_down12 ) ;
  TBCLL pulldown20 ( pull_down20 ) ;
  TBCLL pulldown13 ( pull_down13 ) ;
  TBCLL pulldown21 ( pull_down21 ) ;
  TBCLL pulldown14 ( pull_down14 ) ;
  TBCLL pulldown22 ( pull_down22 ) ;
  TBCLL pulldown30 ( pull_down30 ) ;
  TBCLL pulldown15 ( pull_down15 ) ;
  TBCLL pulldown23 ( pull_down23 ) ;
  TBCLL pulldown31 ( pull_down31 ) ;
  TBCLL pulldown16 ( pull_down16 ) ;
  TBCLL pulldown24 ( pull_down24 ) ;
  TBCLL pulldown32 ( pull_down32 ) ;
  TBCLL pulldown40 ( pull_down40 ) ;
  TBCLL pulldown17 ( pull_down17 ) ;
  TBCLL pulldown25 ( pull_down25 ) ;
  TBCLL pulldown33 ( pull_down33 ) ;
  TBCLL pulldown41 ( pull_down41 ) ;
  TBCLL pulldown18 ( pull_down18 ) ;
  TBCLL pulldown26 ( pull_down26 ) ;
  TBCLL pulldown34 ( pull_down34 ) ;
  TBCLL pulldown42 ( pull_down42 ) ;
  TBCLL pulldown50 ( pull_down50 ) ;
  TBCLL pulldown19 ( pull_down19 ) ;
  TBCLL pulldown27 ( pull_down27 ) ;
  TBCLL pulldown35 ( pull_down35 ) ;
  TBCLL pulldown43 ( pull_down43 ) ;
  TBCLL pulldown51 ( pull_down51 ) ;
  TBCLL pulldown28 ( pull_down28 ) ;
  TBCLL pulldown36 ( pull_down36 ) ;
  TBCLL pulldown44 ( pull_down44 ) ;
  TBCLL pulldown52 ( pull_down52 ) ;
  TBCLL pulldown60 ( pull_down60 ) ;
  TBCLL pulldown29 ( pull_down29 ) ;
  TBCLL pulldown37 ( pull_down37 ) ;
  TBCLL pulldown45 ( pull_down45 ) ;
  TBCLL pulldown53 ( pull_down53 ) ;
  TBCLL pulldown61 ( pull_down61 ) ;
  TBCLL pulldown38 ( pull_down38 ) ;
  TBCLL pulldown46 ( pull_down46 ) ;
  TBCLL pulldown54 ( pull_down54 ) ;
  TBCLL pulldown62 ( pull_down62 ) ;
  TBCLL pulldown70 ( pull_down70 ) ;
  TBCLL pulldown39 ( pull_down39 ) ;
  TBCLL pulldown47 ( pull_down47 ) ;
  TBCLL pulldown55 ( pull_down55 ) ;
  TBCLL pulldown63 ( pull_down63 ) ;
  TBCLL pulldown71 ( pull_down71 ) ;
  TBCLL pulldown48 ( pull_down48 ) ;
  TBCLL pulldown56 ( pull_down56 ) ;
  TBCLL pulldown64 ( pull_down64 ) ;
  TBCLL pulldown72 ( pull_down72 ) ;
  TBCLL pulldown80 ( pull_down80 ) ;
  TBCLL pulldown49 ( pull_down49 ) ;
  TBCLL pulldown57 ( pull_down57 ) ;
  TBCLL pulldown65 ( pull_down65 ) ;
  TBCLL pulldown73 ( pull_down73 ) ;
  TBCLL pulldown81 ( pull_down81 ) ;
  TBCLL pulldown58 ( pull_down58 ) ;
  TBCLL pulldown66 ( pull_down66 ) ;
  TBCLL pulldown74 ( pull_down74 ) ;
  TBCLL pulldown82 ( pull_down82 ) ;
  TBCLL pulldown90 ( pull_down90 ) ;
  TBCLL pulldown59 ( pull_down59 ) ;
  TBCLL pulldown67 ( pull_down67 ) ;
  TBCLL pulldown75 ( pull_down75 ) ;
  TBCLL pulldown83 ( pull_down83 ) ;
  TBCLL pulldown91 ( pull_down91 ) ;
  TBCLL pulldown68 ( pull_down68 ) ;
  TBCLL pulldown76 ( pull_down76 ) ;
  TBCLL pulldown84 ( pull_down84 ) ;
  TBCLL pulldown92 ( pull_down92 ) ;
  TBCLL pulldown69 ( pull_down69 ) ;
  TBCLL pulldown77 ( pull_down77 ) ;
  TBCLL pulldown85 ( pull_down85 ) ;
  TBCLL pulldown93 ( pull_down93 ) ;
  TBCLL pulldown78 ( pull_down78 ) ;
  TBCLL pulldown86 ( pull_down86 ) ;
  TBCLL pulldown94 ( pull_down94 ) ;
  TBCLL pulldown79 ( pull_down79 ) ;
  TBCLL pulldown87 ( pull_down87 ) ;
  TBCLL pulldown95 ( pull_down95 ) ;
  TBCLL pulldown88 ( pull_down88 ) ;
  TBCLL pulldown96 ( pull_down96 ) ;
  TBCLL pulldown89 ( pull_down89 ) ;
  TBCLL pulldown97 ( pull_down97 ) ;
  TBCLL pulldown98 ( pull_down98 ) ;
  TBCLL pulldown99 ( pull_down99 ) ;
  TBCLL pulldown100 ( pull_down100 ) ;
  TBCLL pulldown101 ( pull_down101 ) ;
  TBCLL pulldown102 ( pull_down102 ) ;
  TBCLL pulldown110 ( pull_down110 ) ;
  TBCLL pulldown103 ( pull_down103 ) ;
  TBCLL pulldown111 ( pull_down111 ) ;
  TBCLL pulldown104 ( pull_down104 ) ;
  TBCLL pulldown112 ( pull_down112 ) ;
  TBCLL pulldown120 ( pull_down120 ) ;
  TBCLL pulldown105 ( pull_down105 ) ;
  TBCLL pulldown113 ( pull_down113 ) ;
  TBCLL pulldown106 ( pull_down106 ) ;
  TBCLL pulldown114 ( pull_down114 ) ;
  TBCLL pulldown107 ( pull_down107 ) ;
  TBCLL pulldown115 ( pull_down115 ) ;
  TBCLL pulldown108 ( pull_down108 ) ;
  TBCLL pulldown116 ( pull_down116 ) ;
  TBCLL pulldown109 ( pull_down109 ) ;
  TBCLL pulldown117 ( pull_down117 ) ;
  TBCLL pulldown118 ( pull_down118 ) ;
  TBCLL pulldown119 ( pull_down119 ) ;
  TBCLH pullup0 ( pull_up0 ) ;
  TBCLH pullup1 ( pull_up1 ) ;
  TBCLH pullup2 ( pull_up2 ) ;
  TBCLH pullup3 ( pull_up3 ) ;
  TBCLH pullup4 ( pull_up4 ) ;
  TBCLH pullup5 ( pull_up5 ) ;
  TBCLH pullup6 ( pull_up6 ) ;
  TBCLH pullup7 ( pull_up7 ) ;
  TBCLH pullup8 ( pull_up8 ) ;
  TBCLH pullup9 ( pull_up9 ) ;
  TBCLH pullup10 ( pull_up10 ) ;
  TBCLH pullup11 ( pull_up11 ) ;
  TBCLH pullup12 ( pull_up12 ) ;
  TBCLH pullup20 ( pull_up20 ) ;
  TBCLH pullup13 ( pull_up13 ) ;
  TBCLH pullup21 ( pull_up21 ) ;
  TBCLH pullup14 ( pull_up14 ) ;
  TBCLH pullup22 ( pull_up22 ) ;
  TBCLH pullup30 ( pull_up30 ) ;
  TBCLH pullup15 ( pull_up15 ) ;
  TBCLH pullup23 ( pull_up23 ) ;
  TBCLH pullup31 ( pull_up31 ) ;
  TBCLH pullup16 ( pull_up16 ) ;
  TBCLH pullup24 ( pull_up24 ) ;
  TBCLH pullup32 ( pull_up32 ) ;
  TBCLH pullup40 ( pull_up40 ) ;
  TBCLH pullup17 ( pull_up17 ) ;
  TBCLH pullup25 ( pull_up25 ) ;
  TBCLH pullup33 ( pull_up33 ) ;
  TBCLH pullup41 ( pull_up41 ) ;
  TBCLH pullup18 ( pull_up18 ) ;
  TBCLH pullup26 ( pull_up26 ) ;
  TBCLH pullup34 ( pull_up34 ) ;
  TBCLH pullup42 ( pull_up42 ) ;
  TBCLH pullup50 ( pull_up50 ) ;
  TBCLH pullup19 ( pull_up19 ) ;
  TBCLH pullup27 ( pull_up27 ) ;
  TBCLH pullup35 ( pull_up35 ) ;
  TBCLH pullup43 ( pull_up43 ) ;
  TBCLH pullup51 ( pull_up51 ) ;
  TBCLH pullup28 ( pull_up28 ) ;
  TBCLH pullup36 ( pull_up36 ) ;
  TBCLH pullup44 ( pull_up44 ) ;
  TBCLH pullup52 ( pull_up52 ) ;
  TBCLH pullup60 ( pull_up60 ) ;
  TBCLH pullup29 ( pull_up29 ) ;
  TBCLH pullup37 ( pull_up37 ) ;
  TBCLH pullup45 ( pull_up45 ) ;
  TBCLH pullup53 ( pull_up53 ) ;
  TBCLH pullup61 ( pull_up61 ) ;
  TBCLH pullup38 ( pull_up38 ) ;
  TBCLH pullup46 ( pull_up46 ) ;
  TBCLH pullup54 ( pull_up54 ) ;
  TBCLH pullup62 ( pull_up62 ) ;
  TBCLH pullup70 ( pull_up70 ) ;
  TBCLH pullup39 ( pull_up39 ) ;
  TBCLH pullup47 ( pull_up47 ) ;
  TBCLH pullup55 ( pull_up55 ) ;
  TBCLH pullup63 ( pull_up63 ) ;
  TBCLH pullup71 ( pull_up71 ) ;
  TBCLH pullup48 ( pull_up48 ) ;
  TBCLH pullup56 ( pull_up56 ) ;
  TBCLH pullup64 ( pull_up64 ) ;
  TBCLH pullup72 ( pull_up72 ) ;
  TBCLH pullup49 ( pull_up49 ) ;
  TBCLH pullup57 ( pull_up57 ) ;
  TBCLH pullup65 ( pull_up65 ) ;
  TBCLH pullup73 ( pull_up73 ) ;
  TBCLH pullup58 ( pull_up58 ) ;
  TBCLH pullup66 ( pull_up66 ) ;
  TBCLH pullup74 ( pull_up74 ) ;
  TBCLH pullup59 ( pull_up59 ) ;
  TBCLH pullup67 ( pull_up67 ) ;
  TBCLH pullup75 ( pull_up75 ) ;
  TBCLH pullup68 ( pull_up68 ) ;
  TBCLH pullup76 ( pull_up76 ) ;
  TBCLH pullup69 ( pull_up69 ) ;
  TBCLH pullup77 ( pull_up77 ) ;
  TBCLH pullup78 ( pull_up78 ) ;
  TBCLH pullup79 ( pull_up79 ) ;

  // Refer to /proj/78k0r_3/ss2/_macro/qlk0rcpueva0v3_mf3_v3.10/_library/qlk0rcpueva0v3_101216.hdl
  QLK0RCPUEVA0V3 cpu (
    .PC19 ( PC19 ) ,.PC18 ( PC18 ) ,.PC17 ( PC17 ) ,.PC16 ( PC16 ) ,.PC15 ( PC15 )
     ,.PC14 ( PC14 ) ,.PC13 ( PC13 ) ,.PC12 ( PC12 ) ,.PC11 ( PC11 ) ,.PA19 ( PA19 )
     ,.PC10 ( PC10 ) ,.PA18 ( PA18 ) ,.PC9 ( PC9 ) ,.PC8 ( PC8 ) ,.PC7 ( PC7 )
     ,.PC6 ( PC6 ) ,.PC5 ( PC5 ) ,.PA9 ( PA9 ) ,.PC4 ( PC4 ) ,.PA8 ( PA8 )
     ,.PC3 ( PC3 ) ,.PA7 ( PA7 ) ,.PC2 ( PC2 ) ,.PA6 ( PA6 ) ,.PC1 ( PC1 )
     ,.PA5 ( PA5 ) ,.PC0 ( PC0 ) ,.PA4 ( PA4 ) ,.PA17 ( PA17 ) ,.PA16 ( PA16 )
     ,.PA15 ( PA15 ) ,.PA14 ( PA14 ) ,.PA13 ( PA13 ) ,.PA12 ( PA12 ) ,.PA11 ( PA11 )
     ,.PA10 ( PA10 ) ,.PA3 ( PA3 ) ,.PA2 ( PA2 ) ,.PID31 ( CPUPID31 ) ,.PID23 ( CPUPID23 )
     ,.PID15 ( CPUPID15 ) ,.PID30 ( CPUPID30 ) ,.PID22 ( CPUPID22 ) ,.PID14 ( CPUPID14 )
     ,.PID29 ( CPUPID29 ) ,.PID28 ( CPUPID28 ) ,.PID27 ( CPUPID27 ) ,.PID19 ( CPUPID19 )
     ,.PID26 ( CPUPID26 ) ,.PID18 ( CPUPID18 ) ,.PID25 ( CPUPID25 ) ,.PID17 ( CPUPID17 )
     ,.PID24 ( CPUPID24 ) ,.PID16 ( CPUPID16 ) ,.PID21 ( CPUPID21 ) ,.PID13 ( CPUPID13 )
     ,.PID20 ( CPUPID20 ) ,.PID12 ( CPUPID12 ) ,.CPURD ( CPURD ) ,.PID11 ( CPUPID11 )
     ,.PID10 ( CPUPID10 ) ,.PID9 ( CPUPID9 ) ,.PID8 ( CPUPID8 ) ,.PID7 ( CPUPID7 )
     ,.PID6 ( CPUPID6 ) ,.PID5 ( CPUPID5 ) ,.PID4 ( CPUPID4 ) ,.PID3 ( CPUPID3 )
     ,.MDW9 ( MDW9 ) ,.PID2 ( CPUPID2 ) ,.MDW8 ( MDW8 ) ,.PID1 ( CPUPID1 )
     ,.MDW7 ( MDW7 ) ,.PID0 ( CPUPID0 ) ,.MDW6 ( MDW6 ) ,.MA15 ( MA15 )
     ,.MA14 ( MA14 ) ,.MA13 ( MA13 ) ,.MA12 ( MA12 ) ,.MA11 ( MA11 ) ,.MA10 ( MA10 )
     ,.MA9 ( MA9 ) ,.MA8 ( MA8 ) ,.MA7 ( MA7 ) ,.MA6 ( MA6 ) ,.MA5 ( MA5 )
     ,.MA4 ( MA4 ) ,.MA3 ( MA3 ) ,.MA2 ( MA2 ) ,.MA1 ( MA1 ) ,.MA0 ( MA0 )
     ,.DMAMA15 ( DMAMA15 ) ,.DMAMA14 ( DMAMA14 ) ,.DMAMA13 ( DMAMA13 )
     ,.DMAMA12 ( DMAMA12 ) ,.DMAMA11 ( DMAMA11 ) ,.DMAMA10 ( DMAMA10 )
     ,.DMAMA9 ( DMAMA9 ) ,.FCHRAM ( FCHRAM ) ,.DMAMA8 ( DMAMA8 ) ,.DMAMA7 ( DMAMA7 )
     ,.DMAMA6 ( DMAMA6 ) ,.DMAMA5 ( DMAMA5 ) ,.DMAMA4 ( DMAMA4 ) ,.DMAMA3 ( DMAMA3 )
     ,.DMAMA2 ( DMAMA2 ) ,.DMAMA1 ( DMAMA1 ) ,.DMAMA0 ( DMAMA0 ) ,.DMARQ ( DMARQ )
     ,.DMAACK ( DMAACK ) ,.DMARD ( DMARD ) ,.DMAWR ( DMAWR ) ,.DMAWDOP ( DMAWDOP )
     ,.DMAEN ( DMAEN ) ,.SLMEM ( SLMEM ) ,.SLFLASH ( SLFLASH ) ,.WAITFL2 ( WAITFL2 )
     ,.SLEXM ( SLEXM ) ,.SLBMEM ( SLBMEM ) ,.SLIRAM ( SLIRAM ) ,.HLTST ( HLTST )
     ,.STPST ( STPST ) ,.STBEN ( STBEN ) ,.MDR15 ( MDR15 ) ,.MDR14 ( MDR14 )
     ,.MDR13 ( MDR13 ) ,.MDR12 ( MDR12 ) ,.MDR11 ( MDR11 ) ,.MDR10 ( MDR10 )
     ,.MDR9 ( MDR9 ) ,.MDR8 ( MDR8 ) ,.MDR7 ( MDR7 ) ,.MDR6 ( MDR6 ) ,.MDR5 ( MDR5 )
     ,.MDR4 ( MDR4 ) ,.MDR3 ( MDR3 ) ,.MDR2 ( MDR2 ) ,.MDR1 ( MDR1 ) ,.MDR0 ( MDR0 )
     ,.MDW15 ( MDW15 ) ,.IMDR7 ( IMDR7 ) ,.MDW14 ( MDW14 ) ,.IMDR6 ( IMDR6 )
     ,.MDW13 ( MDW13 ) ,.IMDR5 ( IMDR5 ) ,.MDW12 ( MDW12 ) ,.IMDR4 ( IMDR4 )
     ,.MDW11 ( MDW11 ) ,.IMDR3 ( IMDR3 ) ,.MDW10 ( MDW10 ) ,.IDPOP ( IDPOP )
     ,.IMDR2 ( IMDR2 ) ,.MDW5 ( MDW5 ) ,.MDW4 ( MDW4 ) ,.MDW3 ( MDW3 )
     ,.MDW2 ( MDW2 ) ,.MDW1 ( MDW1 ) ,.MDW0 ( MDW0 ) ,.BITEN7 ( BITEN7 )
     ,.ICEDO1 ( ICEDO1 ) ,.BITEN6 ( BITEN6 ) ,.ICEDO0 ( ICEDO0 ) ,.BITEN5 ( BITEN5 )
     ,.IDADR9 ( IDADR9 ) ,.BITEN4 ( BITEN4 ) ,.IDADR8 ( IDADR8 ) ,.BITEN3 ( BITEN3 )
     ,.IDADR7 ( IDADR7 ) ,.BITEN2 ( BITEN2 ) ,.IDADR6 ( IDADR6 ) ,.BITEN1 ( BITEN1 )
     ,.IDADR5 ( IDADR5 ) ,.BITEN0 ( BITEN0 ) ,.IDADR4 ( IDADR4 ) ,.CPUWR ( CPUWR )
     ,.WDOP ( WDOP ) ,.WDWR ( WDWR ) ,.EXMA3 ( EXMA3 ) ,.FLSPM ( FLSPM )
     ,.EXMA2 ( EXMA2 ) ,.EXMA1 ( EXMA1 ) ,.EXMA0 ( EXMA0 ) ,.VCOUT6 ( VCOUT6 )
     ,.VCOUT5 ( VCOUT5 ) ,.VCOUT4 ( VCOUT4 ) ,.VCOUT3 ( VCOUT3 ) ,.VCOUT2 ( VCOUT2 )
     ,.VCOUT1 ( VCOUT1 ) ,.INTDBG ( INTDBG ) ,.INTNMI ( INTNMI ) ,.INTRQ1 ( INTRQ1 )
     ,.INTRQ3 ( INTRQ3 ) ,.INTRQ2 ( INTRQ2 ) ,.INTRQ0 ( INTRQ0 ) ,.INTACK ( INTACK )
     ,.SKIPEXE ( SKIPEXE ) ,.MONMD ( MONMD ) ,.MONMDSTP ( MONMDSTP ) ,.SOFTBRK ( SOFTBRK )
     ,.BRKMSK ( BRKMSK ) ,.WAITMEM ( BBWAITMEM ) ,.WAITFL ( pull_down7 )
     ,.WAITMOD ( WAITMOD ) ,.WAITEXM ( pull_down6 ) ,.DMAWAIT ( DMAWAIT )
     ,.OCDWAIT ( OCDWAIT ) ,.FLSIZE3 ( FLSIZE3 ) ,.FLSIZE2 ( FLSIZE2 )
     ,.FLSIZE1 ( FLSIZE1 ) ,.FLSIZE0 ( FLSIZE0 ) ,.BFSIZE3 ( BFSIZE3 )
     ,.BFSIZE2 ( BFSIZE2 ) ,.BFSIZE1 ( BFSIZE1 ) ,.BFSIZE0 ( BFSIZE0 )
     ,.RAMSIZE7 ( RAMSIZE7 ) ,.RAMSIZE6 ( RAMSIZE6 ) ,.RAMSIZE5 ( RAMSIZE5 )
     ,.RAMSIZE4 ( RAMSIZE4 ) ,.RAMSIZE3 ( RAMSIZE3 ) ,.RAMSIZE2 ( RAMSIZE2 )
     ,.RAMSIZE1 ( RAMSIZE1 ) ,.RAMSIZE0 ( RAMSIZE0 ) ,.BMSIZE3 ( BMSIZE3 )
     ,.BMSIZE2 ( BMSIZE2 ) ,.BMSIZE1 ( BMSIZE1 ) ,.BMSIZE0 ( BMSIZE0 )
     ,.WAIT2ND7 ( pull_down0 ) ,.WAIT2ND6 ( BBWAIT56 ) ,.WAIT2ND5 ( BBWAIT56 )
     ,.WAIT2ND4 ( pull_down1 ) ,.WAIT2ND3 ( pull_down2 ) ,.WAIT2ND2 ( pull_down3 )
     ,.WAIT2ND1 ( pull_down4 ) ,.WAIT2ND0 ( pull_down5 ) ,.FLREAD ( FLREAD )
     ,.IMDR10 ( IMDR10 ) ,.ICEWAITMEM ( ICEWAITMEM ) ,.SVI ( SVI ) ,.SVVCOUT7 ( SVVCOUT7 )
     ,.SVVCOUT6 ( SVVCOUT6 ) ,.SVVCOUT5 ( SVVCOUT5 ) ,.SVVCOUT4 ( SVVCOUT4 )
     ,.SVVCOUT3 ( SVVCOUT3 ) ,.SVVCOUT2 ( SVVCOUT2 ) ,.SVVCOUT1 ( SVVCOUT1 )
     ,.SVVCOUT0 ( SVVCOUT0 ) ,.SVINTACK ( SVINTACK ) ,.SVMOD ( SVMOD )
     ,.SVMODF ( SVMODF ) ,.ALT1 ( ALT1 ) ,.ALT2 ( ALT2 ) ,.SP15 ( SP15 )
     ,.SP14 ( SP14 ) ,.SP13 ( SP13 ) ,.SP12 ( SP12 ) ,.SP11 ( SP11 ) ,.SP10 ( SP10 )
     ,.SP9 ( SP9 ) ,.SP8 ( SP8 ) ,.SP7 ( SP7 ) ,.SP6 ( SP6 ) ,.SP5 ( SP5 )
     ,.SP4 ( SP4 ) ,.SP3 ( SP3 ) ,.SP2 ( SP2 ) ,.SP1 ( SP1 ) ,.SP0 ( SP0 )
     ,.SPINC ( SPINC ) ,.SPDEC ( SPDEC ) ,.ICECSGREGU ( ICECSGREGU ) ,.ICECSGREGA ( pull_down8 )
     ,.ICEIFA4 ( ICEIFA4 ) ,.GATEAD2 ( MONACTIVE ) ,.ICEIFA3 ( ICEIFA3 )
     ,.GATEAD1 ( OCDMOD ) ,.ICEIFA2 ( ICEIFA2 ) ,.ICEDO31 ( ICEDO31 ) ,.ICEDO23 ( ICEDO23 )
     ,.ICEDO15 ( ICEDO15 ) ,.ICEDO30 ( ICEDO30 ) ,.ICEDO22 ( ICEDO22 )
     ,.ICEDO14 ( ICEDO14 ) ,.ICEDO29 ( ICEDO29 ) ,.ICEDO28 ( ICEDO28 )
     ,.ICEDO27 ( ICEDO27 ) ,.ICEDO19 ( ICEDO19 ) ,.ICEDO26 ( ICEDO26 )
     ,.ICEDO18 ( ICEDO18 ) ,.ICEDO25 ( ICEDO25 ) ,.ICEDO17 ( ICEDO17 )
     ,.ICEDO24 ( ICEDO24 ) ,.ICEDO16 ( ICEDO16 ) ,.ICEDO21 ( ICEDO21 )
     ,.ICEDO13 ( ICEDO13 ) ,.ICEDO20 ( ICEDO20 ) ,.ICEDO12 ( ICEDO12 )
     ,.ICEDO11 ( ICEDO11 ) ,.ICEDO10 ( ICEDO10 ) ,.ICEDO9 ( ICEDO9 ) ,.ICEDO8 ( ICEDO8 )
     ,.ICEDO7 ( ICEDO7 ) ,.ICEDO6 ( ICEDO6 ) ,.ICEDO5 ( ICEDO5 ) ,.ICEDO4 ( ICEDO4 )
     ,.ICEDO3 ( ICEDO3 ) ,.ICEDO2 ( ICEDO2 ) ,.FLREADB3 ( FLREADB3 ) ,.FLREADB2 ( FLREADB2 )
     ,.FLREADB1 ( FLREADB1 ) ,.FLREADB0 ( FLREADB0 ) ,.IMDR15 ( IMDR15 )
     ,.IMDR14 ( IMDR14 ) ,.IMDR13 ( IMDR13 ) ,.IMDR12 ( IMDR12 ) ,.IMDR11 ( IMDR11 )
     ,.IMDR9 ( IMDR9 ) ,.IMDR8 ( IMDR8 ) ,.IMDR1 ( IMDR1 ) ,.IMDR0 ( IMDR0 )
     ,.IDADR31 ( IDADR31 ) ,.IDADR23 ( IDADR23 ) ,.IDADR15 ( IDADR15 )
     ,.IDADR30 ( IDADR30 ) ,.IDADR22 ( IDADR22 ) ,.IDADR14 ( IDADR14 )
     ,.IDADR29 ( IDADR29 ) ,.IDADR28 ( IDADR28 ) ,.IDADR27 ( IDADR27 )
     ,.IDADR19 ( IDADR19 ) ,.IDADR26 ( IDADR26 ) ,.IDADR18 ( IDADR18 )
     ,.IDADR25 ( IDADR25 ) ,.IDADR17 ( IDADR17 ) ,.IDADR24 ( IDADR24 )
     ,.IDADR16 ( IDADR16 ) ,.IDADR21 ( IDADR21 ) ,.IDADR13 ( IDADR13 )
     ,.IDADR20 ( IDADR20 ) ,.IDADR12 ( IDADR12 ) ,.IDADR11 ( IDADR11 )
     ,.IDADR10 ( IDADR10 ) ,.IDADR3 ( IDADR3 ) ,.IDADR2 ( IDADR2 ) ,.IDADR1 ( IDADR1 )
     ,.IDADR0 ( IDADR0 ) ,.STAGEADR1 ( STAGEADR1 ) ,.STAGEADR0 ( STAGEADR0 )
     ,.PREFIX ( PREFIX ) ,.PCWAITF ( PCWAITF ) ,.ICEMSKNMI ( ICEMSKNMI )
     ,.ICEMSKDBG ( ICEMSKDBG ) ,.CPUMASK ( CPUMASK ) ,.CPUMISAL ( CPUMISAL )
     ,.SPREL ( SPREL ) ,.OCDMOD ( OCDMOD ) ,.PSELCPU ( PSELCPU ) ,.PSELBCD ( PSELBCD )
     ,.CPUSTART ( CPUSTART ) ,.BASECKHS ( BASECKHS ) ,.RESB ( RESB ) ,.SCANMODE ( SCANMODE )
     ,.DFSIZE1 ( DFSIZE1 ) ,.DFSIZE0 ( DFSIZE0 ) ,.DFLEN ( DFLEN ) ,.SLDFLASH ( SLDFLASH )
     ,.DRDCLK ( DRDCLK ) ,.WED ( WED ) ,.GOFIRM ( GOFIRM ) ,.GATEAD3 ( CSPDTFLG )
     ,.MONPC19 ( MONPC19 ) ,.MONPC18 ( MONPC18 ) ,.MONPC17 ( MONPC17 )
     ,.MONPC16 ( MONPC16 ) ,.MONPC15 ( MONPC15 ) ,.MONPC14 ( MONPC14 )
     ,.MONPC13 ( MONPC13 ) ,.MONPC12 ( MONPC12 ) ,.MONPC11 ( MONPC11 )
     ,.MONPC10 ( MONPC10 ) ,.MONPC9 ( MONPC9 ) ,.MONPC8 ( MONPC8 ) ,.MONPC7 ( MONPC7 )
     ,.MONPC6 ( MONPC6 ) ,.MONPC5 ( MONPC5 ) ,.MONPC4 ( MONPC4 ) ,.MONPC3 ( MONPC3 )
     ,.MONPC2 ( MONPC2 ) ,.MONPC1 ( MONPC1 ) ,.MONPC0 ( MONPC0 ) ,.MONMA15 ( MONMA15 )
     ,.MONMA14 ( MONMA14 ) ,.MONMA13 ( MONMA13 ) ,.MONMA12 ( MONMA12 )
     ,.MONMA11 ( MONMA11 ) ,.MONMA10 ( MONMA10 ) ,.MONMA9 ( MONMA9 ) ,.MONMA8 ( MONMA8 )
     ,.MONMA7 ( MONMA7 ) ,.MONMA6 ( MONMA6 ) ,.MONMA5 ( MONMA5 ) ,.MONMA4 ( MONMA4 )
     ,.MONMA3 ( MONMA3 ) ,.MONMA2 ( MONMA2 ) ,.MONMA1 ( MONMA1 ) ,.MONMA0 ( MONMA0 )
     ,.MONMDR15 ( MONMDR15 ) ,.MONMDR14 ( MONMDR14 ) ,.MONMDR13 ( MONMDR13 )
     ,.MONMDR12 ( MONMDR12 ) ,.MONMDR11 ( MONMDR11 ) ,.MONMDR10 ( MONMDR10 )
     ,.MONMDR9 ( MONMDR9 ) ,.MONMDR8 ( MONMDR8 ) ,.MONMDR7 ( MONMDR7 )
     ,.MONMDR6 ( MONMDR6 ) ,.MONMDR5 ( MONMDR5 ) ,.MONMDR4 ( MONMDR4 )
     ,.MONMDR3 ( MONMDR3 ) ,.MONMDR2 ( MONMDR2 ) ,.MONMDR1 ( MONMDR1 )
     ,.MONMDR0 ( MONMDR0 ) ,.MONMDW15 ( MONMDW15 ) ,.MONMDW14 ( MONMDW14 )
     ,.MONMDW13 ( MONMDW13 ) ,.MONMDW12 ( MONMDW12 ) ,.MONMDW11 ( MONMDW11 )
     ,.MONMDW10 ( MONMDW10 ) ,.MONMDW9 ( MONMDW9 ) ,.MONMDW8 ( MONMDW8 )
     ,.MONMDW7 ( MONMDW7 ) ,.MONMDW6 ( MONMDW6 ) ,.MONMDW5 ( MONMDW5 )
     ,.MONMDW4 ( MONMDW4 ) ,.MONMDW3 ( MONMDW3 ) ,.MONMDW2 ( MONMDW2 )
     ,.MONMDW1 ( MONMDW1 ) ,.MONMDW0 ( MONMDW0 ) ,.CRCHLTEN ( CRCHLTEN )
    
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_soft/qlk0rint48v2_mf3_v2.10/_library/100722/qlk0rint48v2.hdl
  QLK0RINT48V2 int48 (
    .INTAS02 ( INTAS02 ) ,.INTAS10 ( INTP4 ) ,.INTAS04 ( INTAS04 ) ,.INTAS12 ( INTP5 )
     ,.INTAS20 ( INTSAU01 ) ,.INTAS06 ( INTLVI ) ,.INTAS14 ( INTSAU10 )
     ,.INTAS22 ( INTAS22 ) ,.INTAS30 ( INTTM02 ) ,.INTAS08 ( INTP0 ) ,.INTAS16 ( INTSAU11 )
     ,.INTAS24 ( INTSAU02 ) ,.INTAS32 ( INTTM03 ) ,.INTAS40 ( BBINT2 )
     ,.INTAS0A ( INTP1 ) ,.INTAS0C ( INTP2 ) ,.INTAS1A ( INTDMA0 ) ,.INTAS0E ( INTP3 )
     ,.INTAS1C ( INTDMA1 ) ,.INTAS2A ( INTIIC0 ) ,.INTAS18 ( INTSRE2 )
     ,.INTAS26 ( INTSAU03 ) ,.INTAS34 ( INTAD ) ,.INTAS42 ( INTTM04 ) ,.INTAS50 ( INTAS50 )
     ,.INTAS1E ( INTSAU00 ) ,.INTAS2C ( INTTM00 ) ,.INTAS3A ( INTKR ) ,.INTAS28 ( INTAS28 )
     ,.INTAS36 ( INTRTC ) ,.INTAS44 ( INTTM05 ) ,.INTAS52 ( INTAS52 ) ,.INTAS60 ( BBINT13 )
     ,.INTAS2E ( INTTM01 ) ,.INTAS3C ( BBINT0 ) ,.INTAS4A ( INTAS4A ) ,.INTAS38 ( INTRTCI )
     ,.INTAS46 ( INTTM06 ) ,.INTAS54 ( INTAS54 ) ,.INTAS62 ( INTFL ) ,.INTAS3E ( BBINT1 )
     ,.INTAS4C ( INTAS4C ) ,.INTAS5A ( BBINT11 ) ,.INTAS48 ( INTTM07 )
     ,.INTAS56 ( BBINT9 ) ,.INTAS4E ( INTAS4E ) ,.INTAS5C ( BBINT12 ) ,.INTAS58 ( BBINT10 )
     ,.INTAS5E ( INTMD ) ,.INTS04EN ( pull_up0 ) ,.INTS12EN ( pull_up7 )
     ,.INTS20EN ( pull_up14 ) ,.INTS06EN ( pull_up1 ) ,.INTS14EN ( pull_up8 )
     ,.INTS22EN ( pull_up15 ) ,.INTS30EN ( pull_up22 ) ,.INTS08EN ( pull_up2 )
     ,.INTS16EN ( pull_up9 ) ,.INTS24EN ( pull_up16 ) ,.INTS32EN ( pull_up23 )
     ,.INTS40EN ( pull_up30 ) ,.INTS0AEN ( pull_up3 ) ,.INTS0CEN ( pull_up4 )
     ,.INTS1AEN ( pull_up11 ) ,.INTS0EEN ( pull_up5 ) ,.INTS1CEN ( pull_up12 )
     ,.INTS2AEN ( pull_up19 ) ,.INTS10EN ( pull_up6 ) ,.INTS18EN ( pull_up10 )
     ,.INTS26EN ( pull_up17 ) ,.INTS34EN ( pull_up24 ) ,.INTS42EN ( pull_up31 )
     ,.INTS50EN ( pull_up38 ) ,.INTS1EEN ( pull_up13 ) ,.INTS2CEN ( pull_up20 )
     ,.INTS3AEN ( pull_up27 ) ,.INTS28EN ( pull_up18 ) ,.INTS36EN ( pull_up25 )
     ,.INTS44EN ( pull_up32 ) ,.INTS52EN ( pull_up39 ) ,.INTS60EN ( pull_up46 )
     ,.INTS2EEN ( pull_up21 ) ,.INTS3CEN ( pull_up28 ) ,.INTS4AEN ( pull_up35 )
     ,.INTS38EN ( pull_up26 ) ,.INTS46EN ( pull_up33 ) ,.INTS54EN ( pull_up40 )
     ,.INTS62EN ( pull_up47 ) ,.INTS3EEN ( pull_up29 ) ,.INTS4CEN ( pull_up36 )
     ,.INTS5AEN ( pull_up43 ) ,.INTS48EN ( pull_up34 ) ,.INTS56EN ( pull_up41 )
     ,.INTS4EEN ( pull_up37 ) ,.INTS5CEN ( pull_up44 ) ,.INTS58EN ( pull_up42 )
     ,.INTS5EEN ( pull_up45 ) ,.NMIMODE ( pull_down9 ) ,.INTDBG ( INTDBG )
     ,.INTNMI ( INTNMI ) ,.INTRQ1 ( INTRQ1 ) ,.INTRQ0 ( INTRQ0 ) ,.INTRQ2 ( INTRQ2 )
     ,.INTRQ3 ( INTRQ3 ) ,.INTACK ( INTACK ) ,.VCOUT6 ( VCOUT6 ) ,.VCOUT5 ( VCOUT5 )
     ,.VCOUT4 ( VCOUT4 ) ,.VCOUT3 ( VCOUT3 ) ,.VCOUT2 ( VCOUT2 ) ,.VCOUT1 ( VCOUT1 )
     ,.STBRELE ( STBRELE ) ,.PSELINT1 ( PSELINT1 ) ,.MA4 ( MA4 ) ,.MA3 ( MA3 )
     ,.MA2 ( MA2 ) ,.MA1 ( MA1 ) ,.MA0 ( MA0 ) ,.MDR15 ( MDRINT15 ) ,.MDR14 ( MDRINT14 )
     ,.MDR13 ( MDRINT13 ) ,.MDR12 ( MDRINT12 ) ,.MDR11 ( MDRINT11 ) ,.MDR10 ( MDRINT10 )
     ,.MDR9 ( MDRINT9 ) ,.MDR8 ( MDRINT8 ) ,.MDR7 ( MDRINT7 ) ,.MDR6 ( MDRINT6 )
     ,.MDR5 ( MDRINT5 ) ,.MDR4 ( MDRINT4 ) ,.MDR3 ( MDRINT3 ) ,.MDR2 ( MDRINT2 )
     ,.MDR1 ( MDRINT1 ) ,.MDR0 ( MDRINT0 ) ,.MDW15 ( MDW15 ) ,.MDW14 ( MDW14 )
     ,.MDW13 ( MDW13 ) ,.MDW12 ( MDW12 ) ,.MDW11 ( MDW11 ) ,.MDW10 ( MDW10 )
     ,.MDW9 ( MDW9 ) ,.MDW8 ( MDW8 ) ,.MDW7 ( MDW7 ) ,.MDW6 ( MDW6 ) ,.MDW5 ( MDW5 )
     ,.MDW4 ( MDW4 ) ,.MDW3 ( MDW3 ) ,.MDW2 ( MDW2 ) ,.MDW1 ( MDW1 ) ,.MDW0 ( MDW0 )
     ,.CPURD ( CPURD ) ,.CPUWR ( CPUWR ) ,.WDOP ( WDOP ) ,.BITEN7 ( BITEN7 )
     ,.BITEN6 ( BITEN6 ) ,.BITEN5 ( BITEN5 ) ,.BITEN4 ( BITEN4 ) ,.BITEN3 ( BITEN3 )
     ,.BITEN2 ( BITEN2 ) ,.BITEN1 ( BITEN1 ) ,.BITEN0 ( BITEN0 ) ,.BASECKHS ( BASECKHS )
     ,.RESB ( RESB ) ,.SCANMODE ( SCANMODE ) ,.SCANCLK ( SCANCLK ) ,.PCLKRW ( PCLKRW )
    
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_1.0/_macro/_soft/qlk0rdmac0v1_mf3_v1.20/_library/091210_df2.0/qlk0rdmac0v1.hdl
  QLK0RDMAC0V1 dmac (
    .PSELDMAC ( PSELDMAC ) ,.MA3 ( MA3 ) ,.MA2 ( MA2 ) ,.MA1 ( MA1 ) ,.MA0 ( MA0 )
     ,.MDW15 ( MDW15 ) ,.MDW14 ( MDW14 ) ,.MDW13 ( MDW13 ) ,.MDW12 ( MDW12 )
     ,.MDW11 ( MDW11 ) ,.MDW10 ( MDW10 ) ,.MDW9 ( MDW9 ) ,.MDW8 ( MDW8 )
     ,.MDW7 ( MDW7 ) ,.MDW6 ( MDW6 ) ,.MDW5 ( MDW5 ) ,.MDW4 ( MDW4 ) ,.MDW3 ( MDW3 )
     ,.MDW2 ( MDW2 ) ,.MDW1 ( MDW1 ) ,.MDW0 ( MDW0 ) ,.MDR15 ( MDRDMA15 )
     ,.MDR14 ( MDRDMA14 ) ,.MDR13 ( MDRDMA13 ) ,.MDR12 ( MDRDMA12 ) ,.MDR11 ( MDRDMA11 )
     ,.MDR10 ( MDRDMA10 ) ,.MDR9 ( MDRDMA9 ) ,.MDR8 ( MDRDMA8 ) ,.MDR7 ( MDRDMA7 )
     ,.MDR6 ( MDRDMA6 ) ,.MDR5 ( MDRDMA5 ) ,.MDR4 ( MDRDMA4 ) ,.MDR3 ( MDRDMA3 )
     ,.MDR2 ( MDRDMA2 ) ,.MDR1 ( MDRDMA1 ) ,.MDR0 ( MDRDMA0 ) ,.CPUWR ( CPUWR )
     ,.CPURD ( CPURD ) ,.WDOP ( WDOP ) ,.TRIGER14 ( INTSRO ) ,.TRIGER13 ( BBINT13 )
     ,.TRIGER12 ( pull_down11 ) ,.TRIGER11 ( pull_down10 ) ,.TRIGER10 ( INTSAU11 )
     ,.TRIGER9 ( INTSAU10 ) ,.TRIGER8 ( INTSAU03 ) ,.TRIGER7 ( INTSAU02 )
     ,.TRIGER6 ( INTSAU01 ) ,.TRIGER5 ( INTSAU00 ) ,.TRIGER4 ( INTTM03 )
     ,.TRIGER3 ( INTTM02 ) ,.TRIGER2 ( INTTM01 ) ,.TRIGER1 ( INTTM00 )
     ,.TRIGER0 ( INTAD ) ,.DMARQ ( DMARQ ) ,.DMAACK ( DMAACK ) ,.DMAMA15 ( DMAMA15 )
     ,.DMAMA14 ( DMAMA14 ) ,.DMAMA13 ( DMAMA13 ) ,.DMAMA12 ( DMAMA12 )
     ,.DMAMA11 ( DMAMA11 ) ,.DMAMA10 ( DMAMA10 ) ,.DMAMA9 ( DMAMA9 ) ,.DMAMA8 ( DMAMA8 )
     ,.DMAMA7 ( DMAMA7 ) ,.DMAMA6 ( DMAMA6 ) ,.DMAMA5 ( DMAMA5 ) ,.DMAMA4 ( DMAMA4 )
     ,.DMAMA3 ( DMAMA3 ) ,.DMAMA2 ( DMAMA2 ) ,.DMAMA1 ( DMAMA1 ) ,.DMAMA0 ( DMAMA0 )
     ,.DMARD ( DMARD ) ,.DMAWR ( DMAWR ) ,.DMAWDOP ( DMAWDOP ) ,.INTDMA0 ( INTDMA0 )
     ,.INTDMA1 ( INTDMA1 ) ,.DMAWAIT ( DMAWAIT ) ,.DMAEN ( DMAEN ) ,.DMACK ( BASECK )
     ,.RESB ( RESB ) ,.SVSTOP ( SVSTOP ) ,.SCANMODE ( SCANMODE )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_1.0/_macro/_soft/qlk0rmuldiv1v1_mf3_v1.00/_library/100129/qlk0rmuldiv1v1.hdl
  QLK0RMULDIV1V1 muldiv (
    .CPURD ( CPURD ) ,.CPUWR ( CPUWR ) ,.PSELMD1 ( PSELMD1 ) ,.PSELMD2 ( PSELMD2 )
     ,.MDW15 ( MDW15 ) ,.MDW14 ( MDW14 ) ,.MDW13 ( MDW13 ) ,.MDW12 ( MDW12 )
     ,.MDW11 ( MDW11 ) ,.MDW10 ( MDW10 ) ,.MDW9 ( MDW9 ) ,.MDW8 ( MDW8 )
     ,.MDW7 ( MDW7 ) ,.MDW6 ( MDW6 ) ,.MDW5 ( MDW5 ) ,.MDW4 ( MDW4 ) ,.MDW3 ( MDW3 )
     ,.MDW2 ( MDW2 ) ,.MDW1 ( MDW1 ) ,.MDW0 ( MDW0 ) ,.MDR15 ( MDRMUL15 )
     ,.MDR14 ( MDRMUL14 ) ,.MDR13 ( MDRMUL13 ) ,.MDR12 ( MDRMUL12 ) ,.MDR11 ( MDRMUL11 )
     ,.MDR10 ( MDRMUL10 ) ,.MDR9 ( MDRMUL9 ) ,.MDR8 ( MDRMUL8 ) ,.MDR7 ( MDRMUL7 )
     ,.MDR6 ( MDRMUL6 ) ,.MDR5 ( MDRMUL5 ) ,.MDR4 ( MDRMUL4 ) ,.MDR3 ( MDRMUL3 )
     ,.MDR2 ( MDRMUL2 ) ,.MDR1 ( MDRMUL1 ) ,.MDR0 ( MDRMUL0 ) ,.MA3 ( MA3 )
     ,.MA2 ( MA2 ) ,.MA1 ( MA1 ) ,.MA0 ( MA0 ) ,.BASECK ( BASECK ) ,.RESB ( RESB )
     ,.SVSTOP ( SVSTOP ) ,.INTMD ( INTMD ) ,.SCANMODE ( SCANMODE ) ,.PCLKRW ( PCLKRW )
    
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_soft/qlk0rocd1v1_mf3_v1.10/_library/100719/qlk0rocd1v1.hdl
  QLK0ROCD1V1 ocd (
    .MONMDR15 ( MONMDR15 ) ,.MONMDR14 ( MONMDR14 ) ,.MONMDR13 ( MONMDR13 )
     ,.MONMDR12 ( MONMDR12 ) ,.MONMDR11 ( MONMDR11 ) ,.MONMDR10 ( MONMDR10 )
     ,.MONMDR9 ( MONMDR9 ) ,.MONMDR8 ( MONMDR8 ) ,.MONMDR7 ( MONMDR7 )
     ,.MONMDR6 ( MONMDR6 ) ,.MONMDR5 ( MONMDR5 ) ,.MONMDR4 ( MONMDR4 )
     ,.MONMDR3 ( MONMDR3 ) ,.MONMDR2 ( MONMDR2 ) ,.MONMDR1 ( MONMDR1 )
     ,.MONMDR0 ( MONMDR0 ) ,.MDR15 ( MDROCD15 ) ,.MDR14 ( MDROCD14 ) ,.MDR13 ( MDROCD13 )
     ,.MDR12 ( MDROCD12 ) ,.MDR11 ( MDROCD11 ) ,.MDR10 ( MDROCD10 ) ,.MDR9 ( MDROCD9 )
     ,.MDR8 ( MDROCD8 ) ,.MDR7 ( MDROCD7 ) ,.MDR6 ( MDROCD6 ) ,.MDR5 ( MDROCD5 )
     ,.MDR4 ( MDROCD4 ) ,.MDR3 ( MDROCD3 ) ,.MDR2 ( MDROCD2 ) ,.MDR1 ( MDROCD1 )
     ,.MDR0 ( MDROCD0 ) ,.MDW15 ( MDW15 ) ,.MDW14 ( MDW14 ) ,.MDW13 ( MDW13 )
     ,.MDW12 ( MDW12 ) ,.MDW11 ( MDW11 ) ,.MDW10 ( MDW10 ) ,.MDW9 ( MDW9 )
     ,.MDW8 ( MDW8 ) ,.MDW7 ( MDW7 ) ,.MDW6 ( MDW6 ) ,.MDW5 ( MDW5 ) ,.MDW4 ( MDW4 )
     ,.MDW3 ( MDW3 ) ,.MDW2 ( MDW2 ) ,.MDW1 ( MDW1 ) ,.MDW0 ( MDW0 ) ,.MONMDW15 ( MONMDW15 )
     ,.MONMDW14 ( MONMDW14 ) ,.MONMDW13 ( MONMDW13 ) ,.MONMDW12 ( MONMDW12 )
     ,.MONMDW11 ( MONMDW11 ) ,.MONMDW10 ( MONMDW10 ) ,.MONMDW9 ( MONMDW9 )
     ,.MONMDW8 ( MONMDW8 ) ,.MONMDW7 ( MONMDW7 ) ,.MONMDW6 ( MONMDW6 )
     ,.MONMDW5 ( MONMDW5 ) ,.MONMDW4 ( MONMDW4 ) ,.MONMDW3 ( MONMDW3 )
     ,.MONMDW2 ( MONMDW2 ) ,.MONMDW1 ( MONMDW1 ) ,.MONMDW0 ( MONMDW0 )
     ,.MONPC19 ( MONPC19 ) ,.MONPC18 ( MONPC18 ) ,.MONPC17 ( MONPC17 )
     ,.MONPC16 ( MONPC16 ) ,.MONPC15 ( MONPC15 ) ,.MONPC14 ( MONPC14 )
     ,.MONPC13 ( MONPC13 ) ,.MONPC12 ( MONPC12 ) ,.MONPC11 ( MONPC11 )
     ,.MONPC10 ( MONPC10 ) ,.MONPC9 ( MONPC9 ) ,.MONPC8 ( MONPC8 ) ,.MONPC7 ( MONPC7 )
     ,.MONPC6 ( MONPC6 ) ,.MONPC5 ( MONPC5 ) ,.MONPC4 ( MONPC4 ) ,.MONPC3 ( MONPC3 )
     ,.MONPC2 ( MONPC2 ) ,.MONPC1 ( MONPC1 ) ,.MONPC0 ( MONPC0 ) ,.MONMA15 ( MONMA15 )
     ,.MONMA14 ( MONMA14 ) ,.MONMA13 ( MONMA13 ) ,.MONMA12 ( MONMA12 )
     ,.MONMA11 ( MONMA11 ) ,.MONMA10 ( MONMA10 ) ,.MONMA9 ( MONMA9 ) ,.MONMA8 ( MONMA8 )
     ,.MONMA7 ( MONMA7 ) ,.MONMA6 ( MONMA6 ) ,.MONMA5 ( MONMA5 ) ,.MONMA4 ( MONMA4 )
     ,.MONMA3 ( MONMA3 ) ,.MONMA2 ( MONMA2 ) ,.MONMA1 ( MONMA1 ) ,.MONMA0 ( MONMA0 )
     ,.MA3 ( MA3 ) ,.MA2 ( MA2 ) ,.MA1 ( MA1 ) ,.MA0 ( MA0 ) ,.PRESOCDZ ( PRESOCDZ )
     ,.PCLKOCD ( PCLKOCD ) ,.CPURD ( CPURD ) ,.CPUWR ( CPUWR ) ,.OCDMOD ( OCDMOD )
     ,.MONMD ( MONSVMOD ) ,.INTAS02 ( INTAS02 ) ,.SVSTOP ( SVSTOPICE )
     ,.SVPERI0 ( SVPERI0ICE ) ,.SVPERI1 ( SVPERI1ICE ) ,.OCDRESMK ( OCDRESMK )
     ,.RXOCD ( RXOCD ) ,.TXOCD ( TXOCD ) ,.SOFTBRK ( SOFTBRK ) ,.OPOCDEN ( OPOCDEN )
     ,.PSELOCD1 ( PSELOCD1 ) ,.PSELOCD2 ( PSELOCD2 ) ,.WDOP ( WDOP ) ,.MONMDSTP ( MONMDSTP )
     ,.SPRGMOD ( SPRGMOD ) ,.SLBMEM ( SLBMEM ) ,.SLMEM ( SLMEM ) ,.INTSRO ( INTSRO )
     ,.OCDWAIT ( OCDWAIT ) ,.SCANMODE ( SCANMODE ) ,.SCANCLK ( SCANCLK )
     ,.SYSRESB ( SYSRESB ) ,.OCDASEN ( OCDASEN ) ,.INTACK ( INTACK ) ,.BRKMSK ( BRKMSK )
     ,.SKIPEXE ( SKIPEXE ) ,.FIHOCD ( FIHOCD ) ,.FRQSEL3 ( FRQSEL3 ) ,.TOOLRX ( P11EXINA )
     ,.SLTRXTX ( SLTRXTX ) ,.GOFIRM ( GOFIRM ) ,.REQOCD ( REQOCD )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_soft/qlk0riaw0v1_mf3_v1.00/_library/100324/qlk0riaw0v1.hdl
  QLK0RIAW0V1 iaw (
    .RESB ( RESB ) ,.BASECKHS ( BASECKHS ) ,.SLEXM ( SLEXM ) ,.SLMEM ( SLMEM )
     ,.CPUWR ( CPUWRIAW ) ,.MONPC19 ( MONPC19 ) ,.MONPC18 ( MONPC18 ) ,.MONPC17 ( MONPC17 )
     ,.MONPC16 ( MONPC16 ) ,.MONPC15 ( MONPC15 ) ,.MONPC14 ( MONPC14 )
     ,.MONPC13 ( MONPC13 ) ,.MONPC12 ( MONPC12 ) ,.MONPC11 ( MONPC11 )
     ,.MONPC10 ( MONPC10 ) ,.MONPC9 ( MONPC9 ) ,.MONPC8 ( MONPC8 ) ,.MONPC7 ( MONPC7 )
     ,.MONPC6 ( MONPC6 ) ,.MONPC5 ( MONPC5 ) ,.MONPC4 ( MONPC4 ) ,.MONMA15 ( MONMA15 )
     ,.MONMA14 ( MONMA14 ) ,.MONMA13 ( MONMA13 ) ,.MONMA12 ( MONMA12 )
     ,.MONMA11 ( MONMA11 ) ,.MONMA10 ( MONMA10 ) ,.MONMA9 ( MONMA9 ) ,.MONMA8 ( MONMA8 )
     ,.MONMA7 ( MONMA7 ) ,.EXMA3 ( EXMA3 ) ,.EXMA2 ( EXMA2 ) ,.EXMA1 ( EXMA1 )
     ,.EXMA0 ( EXMA0 ) ,.SVSTOP ( SVSTOPIAW ) ,.SCANMODE ( SCANMODE ) ,.IAWRES ( IAWRES )
     ,.FLSIZE3 ( FLSIZE3 ) ,.FLSIZE2 ( FLSIZE2 ) ,.FLSIZE1 ( FLSIZE1 )
     ,.FLSIZE0 ( FLSIZE0 ) ,.RAMSIZE7 ( RAMSIZE7 ) ,.RAMSIZE6 ( RAMSIZE6 )
     ,.RAMSIZE5 ( RAMSIZE5 ) ,.RAMSIZE4 ( RAMSIZE4 ) ,.RAMSIZE3 ( RAMSIZE3 )
     ,.RAMSIZE2 ( RAMSIZE2 ) ,.RAMSIZE1 ( RAMSIZE1 ) ,.RAMSIZE0 ( RAMSIZE0 )
     ,.IAWEN ( IAWEN ) ,.OPWDEN ( OPWDEN ) ,.GDRAM1 ( GDRAM1 ) ,.GDRAM0 ( GDRAM0 )
     ,.GDRAMWR ( GDRAMWR ) ,.MONACTIVE ( MONACTIVE )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_soft/qlk0rcsc1v2_mf3_v2.00/_library/100903/qlk0rcsc1v2.hdl
  QLK0RCSC1V2 csc (
    .PSEL3 ( PSELCSC3 ) ,.PSEL2 ( PSELCSC2 ) ,.PSEL1 ( PSELCSC1 ) ,.PADDR2 ( PADDR2 )
     ,.PADDR1 ( PADDR1 ) ,.GOFIRM ( GOFIRM ) ,.PADDR0 ( PADDR0 ) ,.PENABLE ( PENABLE )
     ,.PWRITE ( PWRITE ) ,.PWDATA15 ( MDW15 ) ,.PWDATA14 ( MDW14 ) ,.PWDATA13 ( MDW13 )
     ,.PWDATA12 ( MDW12 ) ,.PWDATA11 ( MDW11 ) ,.PWDATA10 ( MDW10 ) ,.PWDATA9 ( MDW9 )
     ,.PWDATA8 ( MDW8 ) ,.PWDATA7 ( MDW7 ) ,.OPTIDDQ ( OPTIDDQ ) ,.PWDATA6 ( MDW6 )
     ,.PWDATA5 ( MDW5 ) ,.PWDATA4 ( MDW4 ) ,.PWDATA3 ( MDW3 ) ,.PWDATA2 ( MDW2 )
     ,.PWDATA1 ( MDW1 ) ,.OPLVIS1 ( OPLVIS1 ) ,.PWDATA0 ( MDW0 ) ,.OPLVIS0 ( OPLVIS0 )
     ,.OSCOUTM ( OSCOUTM ) ,.OSCOUTS ( OSCOUTS ) ,.R32MOUT ( R32MOUT )
     ,.R15KOUT ( R15KOUT ) ,.EXCLK1 ( EXCLK1 ) ,.SVSTOP ( SVSTOP ) ,.STPST ( STPST )
     ,.HLTST ( HLTST ) ,.STBRELE ( STBRELEICE ) ,.NVMRCEND ( NVMRCEND )
     ,.TESSCAN3 ( TESSCAN3 ) ,.TESSCAN4 ( TESSCAN4 ) ,.OPWDEN ( OPWDEN )
     ,.OPWDSTBY ( OPWDSTBY ) ,.DMAEN ( DMAEN ) ,.OCDMOD ( OCDMOD ) ,.SPRGMOD ( SPRGMOD )
     ,.TESTMOD ( TESTMOD ) ,.PRSCLK8 ( PRSCLK8 ) ,.PTESINST ( PTESINST )
     ,.TESUSR ( TESUSR ) ,.TESDBT ( TESDBT ) ,.PRES1Z ( PRES1Z ) ,.OPTEXCCK ( OPTEXCCK )
     ,.SCANMODE ( SCANMODE ) ,.SCANEN ( SCANEN ) ,.SCANCLK ( SCANCLK )
     ,.SCANRESZ ( SCANRESZ ) ,.POCREL ( POCREL ) ,.RESETB ( RESETB ) ,.POCRELNF ( POCRELNF )
     ,.RESETINBNF ( RESETINBNF ) ,.LVIOUTZNF ( LVIOUTZNF ) ,.WDTRES ( WDTRES )
     ,.SOFTBRK ( PSEUDOON1 ) ,.OCDRESMK ( OCDRESMK ) ,.PRDATA15 ( PRDCSC15 )
     ,.PRDATA14 ( PRDCSC14 ) ,.PRDATA13 ( PRDCSC13 ) ,.PRDATA12 ( PRDCSC12 )
     ,.PRDATA11 ( PRDCSC11 ) ,.PRDATA10 ( PRDCSC10 ) ,.PRDATA9 ( PRDCSC9 )
     ,.PRDATA8 ( PRDCSC8 ) ,.PRDATA7 ( PRDCSC7 ) ,.PRDATA6 ( PRDCSC6 )
     ,.PRDATA5 ( PRDCSC5 ) ,.PRDATA4 ( PRDCSC4 ) ,.PRDATA3 ( PRDCSC3 )
     ,.PRDATA2 ( PRDCSC2 ) ,.PRDATA1 ( PRDCSC1 ) ,.PRDATA0 ( PRDCSC0 )
     ,.BASECK ( BASECK ) ,.BASECKHS ( BASECKHS ) ,.PCLKOCD ( PCLKOCD )
     ,.PCLK7 ( PCLKRTC ) ,.PCLK6 ( PCLK6 ) ,.PCLK5 ( PCLKADC ) ,.PCLK4 ( PCLKIIC )
     ,.PCLK3 ( PCLKSAU1 ) ,.PCLK2 ( PCLKSAU0 ) ,.PCLK1 ( PCLK1 ) ,.PCLK0 ( PCLKTAU0 )
     ,.RESB ( RESB ) ,.NSRESB ( NSRESB ) ,.PRESOCDZ ( PRESOCDZ ) ,.PRESWDTZ ( PRESWDTZ )
     ,.PRES7Z ( PRESRTCZ ) ,.PRES6Z ( PRES6Z ) ,.PRES5Z ( PRESADCZ ) ,.PRES4Z ( PRESIICZ )
     ,.PRES3Z ( PRESSAU1Z ) ,.PRES2Z ( PRESSAU0Z ) ,.PRES0Z ( PRESTAU0Z )
     ,.RESSTP ( RESSTP ) ,.CPUSTART ( CPUSTART ) ,.RESSQSTA ( RESSQSTA )
     ,.FSTPST ( FSTPST ) ,.FHLTST ( FHLTST ) ,.PSUBMODE ( PSUBMODE ) ,.OSCSEL ( OSCSEL )
     ,.MSTOP ( MSTOP ) ,.EXCLK ( EXCLK ) ,.AMPH ( AMPH ) ,.OSCSELS ( OSCSELS )
     ,.XTSTOP ( XTSTOP ) ,.EXCLKS ( EXCLKS ) ,.AMPHS0 ( AMPHS0 ) ,.R32MSTP ( R32MSTP )
     ,.R15KSTPZ ( R15KSTPZ ) ,.REGLC ( REGLC ) ,.REGLV ( REGLV ) ,.OREGSTP ( OREGSTP )
     ,.SYSRESB ( SYSRESB ) ,.LVIEN ( LVIEN ) ,.LVIS2 ( LVIS2 ) ,.LVIS3 ( LVIS3 )
     ,.LVIS1 ( LVIS1 ) ,.LVIS0 ( LVIS0 ) ,.INTLVI ( INTLVI ) ,.TPOCREL ( TPOCREL )
     ,.TLVIF ( TLVIF ) ,.FMAIN ( FMAIN ) ,.PSTN ( PSTN ) ,.AMPHS1 ( AMPHS1 )
     ,.XTWKUP ( XTWKUP ) ,.FCLKRT ( FCLKRT ) ,.SRESREQ ( SRESREQ ) ,.ICECK60M ( ICECK60M )
     ,.ICEMKWDT ( ICEMKWDT ) ,.ICEMKLVI ( ICEMKLVI ) ,.ICEMKSRQ ( ICEMKSRQ )
     ,.TSELOREG ( TSELOREG ) ,.TSELIRES ( TSELIRES ) ,.TTEMP ( TTEMP )
     ,.LOSCTEST ( LOSCTEST ) ,.TSTN ( TSTN ) ,.TFLSTOPC ( TFLSTOPC ) ,.TFLSTOPD ( TFLSTOPD )
     ,.PER07 ( PER07 ) ,.PER06 ( PER06 ) ,.PER05 ( PER05 ) ,.PER04 ( PER04 )
     ,.PER03 ( PER03 ) ,.PER02 ( PER02 ) ,.PER01 ( PER01 ) ,.PER00 ( PER00 )
     ,.STPBCKBT ( STPBCKBT ) ,.CIBRESRQ ( CIBRESRQICE ) ,.OCDASEN ( OCDASEN )
     ,.BBCKSELR ( BBCKSELR ) ,.BBCKSELM ( BBCKSELM ) ,.PCLKRW ( PCLKRW )
     ,.PRSCLK1 ( PRSCLK1 ) ,.PRSCLK2 ( PRSCLK2 ) ,.PRSCLK3 ( PRSCLK3 )
     ,.PRSCLK4 ( PRSCLK4 ) ,.PRSCLK5 ( PRSCLK5 ) ,.PRSCLK6 ( PRSCLK6 )
     ,.PRSCLK7 ( PRSCLK7 ) ,.PRSCLK9 ( PRSCLK9 ) ,.PRSCLK10 ( PRSCLK10 )
     ,.PRSCLK11 ( PRSCLK11 ) ,.PRSCLK12 ( PRSCLK12 ) ,.PRSCLK13 ( PRSCLK13 )
     ,.PRSCLK14 ( PRSCLK14 ) ,.PRSCLK15 ( PRSCLK15 ) ,.RT0LPM ( RT0LPM )
     ,.SVPERI0 ( SVPERI0 ) ,.SVPERI1 ( SVPERI1 ) ,.TMDENCLK ( TMDENCLK )
     ,.FRQSEL4 ( FRQSEL4 ) ,.FRQSEL3 ( FRQSEL3 ) ,.FRQSEL2 ( FRQSEL2 )
     ,.FRQSEL1 ( FRQSEL1 ) ,.FRQSEL0 ( FRQSEL0 ) ,.RDSETUP ( RDSETUP )
     ,.BBCLKR ( BBCLKR ) ,.BBCLKM ( BBCLKM ) ,.INCDECMD ( INCDECMD ) ,.CRCHLTEN ( CRCHLTEN )
     ,.REQPCLKSA ( REQPCLKSAU0 ) ,.REQPCLKAD ( REQPCLKAD ) ,.BBREQPCLK ( BBREQPCLK )
     ,.OPTBCT ( OPTBCT ) ,.REQFL ( REQFL ) ,.REQOCD ( REQOCD ) ,.INTRCLK ( INTRCLK )
     ,.WDTTESCK ( WDTTESCK ) ,.CKSEL ( CKSEL ) ,.CPUCLKEN ( CPUCLKEN )
     ,.RTCCLKEN ( RTCCLKEN ) ,.RPERR ( RPERR ) ,.BBMODE ( BBMODE ) ,.PCLKTST ( PCLKTST )
     ,.IAWRES ( PSEUDOON10 ) ,.SBRFONLY ( SBRFONLY ) ,.FSUB ( FSUB ) ,.STDWAIT ( STDWAIT )
     ,.HISPEED ( HISPEED ) ,.HIOMSK ( HIOMSK ) ,.RLOWSPY ( RLOWSPY ) ,.PAENB ( PAENB )
     ,.OPVPOC2 ( OPVPOC2 ) ,.OPVPOC1 ( OPVPOC1 ) ,.OPVPOC0 ( OPVPOC0 )
     ,.OPLVIMDS1 ( OPLVIMDS1 ) ,.OPLVIMDS0 ( OPLVIMDS0 ) ,.OPBOEN ( OPBOEN )
     ,.LVITEST ( LVITEST ) ,.LVITSEL ( LVITSEL ) ,.PCLKFCB ( PCLKFCB )
     ,.FLROACT ( FLROACT ) ,.FLSPM ( FLSPM ) ,.EEEMD ( EEEMD ) ,.WDEN ( WDEN )
     ,.MCM0 ( MCM0 ) ,.RSTS ( RSTS ) ,.REQR32M ( REQR32M ) ,.VSETEND ( VSETEND )
     ,.BBRPERR ( BBRPERR ) ,.TSELBGR ( TSELBGR ) ,.BBCKSTR ( BBCKSTR )
     ,.PSYSRESB ( PSYSRESB ) ,.BBREGCTL ( BBREGCTL ) ,.BBHIOON ( BBHIOON )
     ,.BBCKSTM ( BBCKSTM ) ,.GOFIRMR ( GOFIRMR ) ,.AMPSEL ( AMPSEL ) ,.FMXST ( FMXST )
     ,.SUBCKST ( SUBCKST ) ,.BCKHSEN ( BCKHSEN ) ,.TRMRD1 ( TRMRD1 )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_1.0/_macro/_soft/qlk0rpclbuz1v1_mf3_v1.00/_library/100210/qlk0rpclbuz1v1.hdl
  QLK0RPCLBUZ1V1 pclbuz (
    .PWDATA15 ( MDW15 ) ,.PWDATA11 ( MDW11 ) ,.PWDATA10 ( MDW10 ) ,.PWDATA9 ( MDW9 )
     ,.PWDATA8 ( MDW8 ) ,.PWDATA7 ( MDW7 ) ,.PWDATA3 ( MDW3 ) ,.PWDATA2 ( MDW2 )
     ,.PWDATA1 ( MDW1 ) ,.PWDATA0 ( MDW0 ) ,.PRDATA15 ( PRDPCL15 ) ,.PRDATA11 ( PRDPCL11 )
     ,.PRDATA10 ( PRDPCL10 ) ,.PRDATA9 ( PRDPCL9 ) ,.PRDATA8 ( PRDPCL8 )
     ,.PRDATA7 ( PRDPCL7 ) ,.PRDATA3 ( PRDPCL3 ) ,.PRDATA2 ( PRDPCL2 )
     ,.PRDATA1 ( PRDPCL1 ) ,.PRDATA0 ( PRDPCL0 ) ,.PADDR0 ( PADDR0 ) ,.PSEL ( PSELPCL )
     ,.PENABLE ( PENABLE ) ,.PWRITE ( PWRITE ) ,.PCLKRW ( PCLKRW ) ,.RESETB ( RESETB )
     ,.RESB ( RESB ) ,.RESSTP ( RESSTP ) ,.FMAIN ( FMAIN ) ,.SCANMODE ( SCANMODE )
     ,.SCANCLK ( SCANCLK ) ,.SCANRESZ ( SCANRESZ ) ,.PCLBUZ0 ( PCLBUZ0 )
     ,.PCLBUZ1 ( PCLBUZ1 ) ,.FSUB ( FSUB )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/_ice/_macro/_sss/cibc/100910/qlk0rcibcevam3sf1v1.hdl
  QLK0RCIBCM3SF1V1 cibc (
    .PENABLE ( PENABLE ) ,.PWRITE ( PWRITE ) ,.PSEL1 ( PSELCIBC ) ,.PADDR3 ( PADDR3 )
     ,.PADDR2 ( PADDR2 ) ,.PADDR1 ( PADDR1 ) ,.PADDR0 ( PADDR0 ) ,.PWDATA15 ( MDW15 )
     ,.PWDATA14 ( MDW14 ) ,.PWDATA13 ( MDW13 ) ,.PWDATA12 ( MDW12 ) ,.PWDATA11 ( MDW11 )
     ,.PWDATA10 ( MDW10 ) ,.PWDATA9 ( MDW9 ) ,.OPWDCS1 ( OPWDCS1 ) ,.PWDATA8 ( MDW8 )
     ,.OPWDCS0 ( OPWDCS0 ) ,.PWDATA7 ( MDW7 ) ,.PWDATA6 ( MDW6 ) ,.PWDATA5 ( MDW5 )
     ,.PWDATA4 ( MDW4 ) ,.PWDATA3 ( MDW3 ) ,.PWDATA2 ( MDW2 ) ,.PWDATA1 ( MDW1 )
     ,.OPLVIS1 ( OPLVIS1 ) ,.PWDATA0 ( MDW0 ) ,.OPLVIS0 ( OPLVIS0 ) ,.PRDATA15 ( PRDCIC15 )
     ,.PRDATA14 ( PRDCIC14 ) ,.PRDATA13 ( PRDCIC13 ) ,.PRDATA12 ( PRDCIC12 )
     ,.PRDATA11 ( PRDCIC11 ) ,.PRDATA10 ( PRDCIC10 ) ,.PRDATA9 ( PRDCIC9 )
     ,.PRDATA8 ( PRDCIC8 ) ,.PRDATA7 ( PRDCIC7 ) ,.PRDATA6 ( PRDCIC6 )
     ,.PRDATA5 ( PRDCIC5 ) ,.PRDATA4 ( PRDCIC4 ) ,.PRDATA3 ( PRDCIC3 )
     ,.PRDATA2 ( PRDCIC2 ) ,.PRDATA1 ( PRDCIC1 ) ,.PRDATA0 ( PRDCIC0 )
     ,.BASECKHS ( BASECKHS ) ,.SYSRESB ( SYSRESB ) ,.RESETB ( RESETB )
     ,.NSRESB ( NSRESB ) ,.PA19 ( PA19 ) ,.PA18 ( PA18 ) ,.CEPR ( CEPR )
     ,.PA17 ( PA17 ) ,.PA16 ( PA16 ) ,.PA15 ( PA15 ) ,.PA14 ( PA14 ) ,.PA13 ( PA13 )
     ,.PA12 ( PA12 ) ,.PA11 ( PA11 ) ,.PA10 ( PA10 ) ,.PA9 ( PA9 ) ,.PA8 ( PA8 )
     ,.PA7 ( PA7 ) ,.PA6 ( PA6 ) ,.PA5 ( PA5 ) ,.PA4 ( PA4 ) ,.PA3 ( PA3 )
     ,.PA2 ( PA2 ) ,.SLFLASH ( SLFLASH ) ,.PID31 ( PID31 ) ,.PID23 ( PID23 )
     ,.PID15 ( PID15 ) ,.RO031 ( RO031 ) ,.RO023 ( RO023 ) ,.RO015 ( RO015 )
     ,.RO111 ( RO111 ) ,.PID30 ( PID30 ) ,.PID22 ( PID22 ) ,.PID14 ( PID14 )
     ,.RO030 ( RO030 ) ,.RO022 ( RO022 ) ,.RO014 ( RO014 ) ,.RO110 ( RO110 )
     ,.PID29 ( PID29 ) ,.RO037 ( RO037 ) ,.RO029 ( RO029 ) ,.RO133 ( RO133 )
     ,.RO125 ( RO125 ) ,.RO117 ( RO117 ) ,.PID28 ( PID28 ) ,.RO036 ( RO036 )
     ,.RO028 ( RO028 ) ,.RO132 ( RO132 ) ,.RO124 ( RO124 ) ,.RO116 ( RO116 )
     ,.PID27 ( PID27 ) ,.PID19 ( PID19 ) ,.RO035 ( RO035 ) ,.RO027 ( RO027 )
     ,.RO019 ( RO019 ) ,.RO131 ( RO131 ) ,.RO123 ( RO123 ) ,.RO115 ( RO115 )
     ,.PID26 ( PID26 ) ,.PID18 ( PID18 ) ,.RO034 ( RO034 ) ,.RO026 ( RO026 )
     ,.RO018 ( RO018 ) ,.RO130 ( RO130 ) ,.RO122 ( RO122 ) ,.RO114 ( RO114 )
     ,.PID25 ( PID25 ) ,.PID17 ( PID17 ) ,.RO033 ( RO033 ) ,.RO025 ( RO025 )
     ,.RO017 ( RO017 ) ,.RO121 ( RO121 ) ,.RO113 ( RO113 ) ,.PID24 ( PID24 )
     ,.PID16 ( PID16 ) ,.RO032 ( RO032 ) ,.RO024 ( RO024 ) ,.RO016 ( RO016 )
     ,.RO120 ( RO120 ) ,.RO112 ( RO112 ) ,.PID21 ( PID21 ) ,.PID13 ( PID13 )
     ,.RO021 ( RO021 ) ,.RO013 ( RO013 ) ,.PID20 ( PID20 ) ,.PID12 ( PID12 )
     ,.RO020 ( RO020 ) ,.RO012 ( RO012 ) ,.PID11 ( PID11 ) ,.RO011 ( RO011 )
     ,.PID10 ( PID10 ) ,.RO010 ( RO010 ) ,.PID9 ( PID9 ) ,.RO09 ( RO09 )
     ,.RO17 ( RO17 ) ,.PID8 ( PID8 ) ,.RO08 ( RO08 ) ,.RO16 ( RO16 ) ,.EXER ( EXER )
     ,.PID7 ( PID7 ) ,.RO07 ( RO07 ) ,.RO15 ( RO15 ) ,.PID6 ( PID6 ) ,.RO06 ( RO06 )
     ,.RO14 ( RO14 ) ,.PID5 ( PID5 ) ,.RO05 ( RO05 ) ,.RO13 ( RO13 ) ,.PID4 ( PID4 )
     ,.RO04 ( RO04 ) ,.RO12 ( RO12 ) ,.PID3 ( PID3 ) ,.RO03 ( RO03 ) ,.RO11 ( RO11 )
     ,.PID2 ( PID2 ) ,.RO02 ( RO02 ) ,.RO10 ( RO10 ) ,.PID1 ( PID1 ) ,.RO01 ( RO01 )
     ,.PID0 ( PID0 ) ,.RO00 ( RO00 ) ,.FHLTST ( FHLTST ) ,.FSTPST ( FSTPST )
     ,.PSUBMODE ( PSUBMODE ) ,.FRSEL4 ( FRSEL4 ) ,.FRSEL3 ( FRSEL3 ) ,.FRSEL2 ( FRSEL2 )
     ,.FLSTOP ( FLSTOP ) ,.FRSEL1 ( FRSEL1 ) ,.FRSEL0 ( FRSEL0 ) ,.OPLVIMDS1 ( OPLVIMDS1 )
     ,.OPLVIMDS0 ( OPLVIMDS0 ) ,.OPVPOC2 ( OPVPOC2 ) ,.OPVPOC1 ( OPVPOC1 )
     ,.OPVPOC0 ( OPVPOC0 ) ,.PORTSELB ( PORTSELB ) ,.OPWDCS2 ( OPWDCS2 )
     ,.OPWDEN ( OPWDEN ) ,.OPWDSTBY ( OPWDSTBY ) ,.OPWDWS1 ( OPWDWS1 )
     ,.OPWDWS0 ( OPWDWS0 ) ,.TMBTSEL ( ICETMBTSEL ) ,.OPWDINT ( OPWDINT )
     ,.OPOCDEN ( OPOCDEN ) ,.C3HFF ( C3HFF ) ,.SELIN1 ( SELIN1 ) ,.AF19 ( AF19 )
     ,.AF18 ( AF18 ) ,.AF17 ( AF17 ) ,.AF16 ( AF16 ) ,.AF15 ( AF15 ) ,.AF14 ( AF14 )
     ,.AF13 ( AF13 ) ,.AF12 ( AF12 ) ,.AF11 ( AF11 ) ,.AF10 ( AF10 ) ,.AF9 ( AF9 )
     ,.AF8 ( AF8 ) ,.AF7 ( AF7 ) ,.CE1 ( CE1 ) ,.AF6 ( AF6 ) ,.CE0 ( CE0 )
     ,.AF5 ( AF5 ) ,.AF4 ( AF4 ) ,.AF3 ( AF3 ) ,.AF2 ( AF2 ) ,.FLRO37 ( FLRO37 )
     ,.FLRO29 ( FLRO29 ) ,.FLRO36 ( FLRO36 ) ,.FLRO28 ( FLRO28 ) ,.FLRO35 ( FLRO35 )
     ,.FLRO27 ( FLRO27 ) ,.FLRO19 ( FLRO19 ) ,.FLRO34 ( FLRO34 ) ,.FLRO26 ( FLRO26 )
     ,.FLRO18 ( FLRO18 ) ,.FLRO33 ( FLRO33 ) ,.FLRO25 ( FLRO25 ) ,.FLRO17 ( FLRO17 )
     ,.FLRO32 ( FLRO32 ) ,.FLRO24 ( FLRO24 ) ,.FLRO16 ( FLRO16 ) ,.FLRO31 ( FLRO31 )
     ,.FLRO23 ( FLRO23 ) ,.FLRO15 ( FLRO15 ) ,.FLRO30 ( FLRO30 ) ,.FLRO22 ( FLRO22 )
     ,.FLRO14 ( FLRO14 ) ,.FLRO21 ( FLRO21 ) ,.FLRO13 ( FLRO13 ) ,.FLRO20 ( FLRO20 )
     ,.FLRO12 ( FLRO12 ) ,.FLRO11 ( FLRO11 ) ,.FLRO10 ( FLRO10 ) ,.FLRO9 ( FLRO9 )
     ,.FLRO8 ( FLRO8 ) ,.FLRO7 ( FLRO7 ) ,.FLRO6 ( FLRO6 ) ,.FLRO5 ( FLRO5 )
     ,.FLRO4 ( FLRO4 ) ,.FLRO3 ( FLRO3 ) ,.FLRO2 ( FLRO2 ) ,.FLRO1 ( FLRO1 )
     ,.FLRO0 ( FLRO0 ) ,.FLSPM ( FLSPM ) ,.RO137 ( RO137 ) ,.RO129 ( RO129 )
     ,.EXCH ( EXCH ) ,.PEXA ( PEXA ) ,.TID9 ( TID9 ) ,.SACEEN ( SACEEN )
     ,.RESSQSTA ( RESSQSTA ) ,.PRDSELEN ( PRDSELEN ) ,.OSCOUTEN ( OSCOUTEN )
     ,.EXCHEN ( EXCHEN ) ,.SECEN ( SECEN ) ,.FSWEN ( FSWEN ) ,.TID20 ( TID20 )
     ,.TID12 ( TID12 ) ,.FSWS2 ( FSWS2 ) ,.NVMRCEND ( NVMRCEND ) ,.TRMCP017 ( TRMCP017 )
     ,.TRMCP113 ( TRMCP113 ) ,.TRMCP016 ( TRMCP016 ) ,.TRMCP112 ( TRMCP112 )
     ,.TRMCP015 ( TRMCP015 ) ,.TRMCP111 ( TRMCP111 ) ,.TRMCP014 ( TRMCP014 )
     ,.TRMCP110 ( TRMCP110 ) ,.TRMCP013 ( TRMCP013 ) ,.TRMCP012 ( TRMCP012 )
     ,.TRMCP011 ( TRMCP011 ) ,.TRMCP010 ( TRMCP010 ) ,.TRMCP09 ( TRMCP09 )
     ,.TRMCP08 ( TRMCP08 ) ,.TRMCP07 ( TRMCP07 ) ,.TRMCP06 ( TRMCP06 )
     ,.TRMCP05 ( TRMCP05 ) ,.TRMCP04 ( TRMCP04 ) ,.TRMCP03 ( TRMCP03 )
     ,.TRMCP02 ( TRMCP02 ) ,.TRMCP01 ( TRMCP01 ) ,.TRMCP00 ( TRMCP00 )
     ,.TRMCP114 ( TRMCP114 ) ,.DTRMCP014 ( DTRMCP014 ) ,.DTRMCP013 ( DTRMCP013 )
     ,.DTRMCP012 ( DTRMCP012 ) ,.DTRMCP011 ( DTRMCP011 ) ,.DTRMCP010 ( DTRMCP010 )
     ,.RTRMCP020 ( RTRMCP020 ) ,.RTRMCP019 ( RTRMCP019 ) ,.RTRMCP018 ( RTRMCP018 )
     ,.RTRMCP017 ( RTRMCP017 ) ,.RTRMCP016 ( RTRMCP016 ) ,.RTRMCP015 ( RTRMCP015 )
     ,.A19 ( A19 ) ,.A18 ( A18 ) ,.A17 ( A17 ) ,.A16 ( A16 ) ,.A15 ( A15 )
     ,.A14 ( A14 ) ,.A13 ( A13 ) ,.A12 ( A12 ) ,.A11 ( A11 ) ,.A10 ( A10 )
     ,.A9 ( A9 ) ,.A8 ( A8 ) ,.A7 ( A7 ) ,.A6 ( A6 ) ,.A5 ( A5 ) ,.A4 ( A4 )
     ,.A3 ( A3 ) ,.A2 ( A2 ) ,.RO136 ( RO136 ) ,.RO128 ( RO128 ) ,.RO135 ( RO135 )
     ,.RO127 ( RO127 ) ,.RO119 ( RO119 ) ,.RO134 ( RO134 ) ,.RO126 ( RO126 )
     ,.RO118 ( RO118 ) ,.RO19 ( RO19 ) ,.RO18 ( RO18 ) ,.EXA ( EXA ) ,.TA3 ( TA3 )
     ,.BFA ( BFA ) ,.CLKSEL1 ( CLKSEL1 ) ,.SRCUT ( SRCUT ) ,.SUB ( SUB )
     ,.HISPEED ( HISPEED ) ,.TID31 ( TID31 ) ,.TID23 ( TID23 ) ,.TID15 ( TID15 )
     ,.FSWS5 ( FSWS5 ) ,.TID30 ( TID30 ) ,.TID22 ( TID22 ) ,.TID14 ( TID14 )
     ,.FSWS4 ( FSWS4 ) ,.TID29 ( TID29 ) ,.TID28 ( TID28 ) ,.TID27 ( TID27 )
     ,.TID19 ( TID19 ) ,.FSWS9 ( FSWS9 ) ,.TID26 ( TID26 ) ,.TID18 ( TID18 )
     ,.FSWS8 ( FSWS8 ) ,.TID25 ( TID25 ) ,.TID17 ( TID17 ) ,.FSWS7 ( FSWS7 )
     ,.TID24 ( TID24 ) ,.TID16 ( TID16 ) ,.FSWS6 ( FSWS6 ) ,.TID21 ( TID21 )
     ,.TID13 ( TID13 ) ,.FSWS3 ( FSWS3 ) ,.TID11 ( TID11 ) ,.FSWS1 ( FSWS1 )
     ,.TID10 ( TID10 ) ,.FSWS0 ( FSWS0 ) ,.TID8 ( TID8 ) ,.TID7 ( TID7 )
     ,.TID6 ( TID6 ) ,.TID5 ( TID5 ) ,.TID4 ( TID4 ) ,.TID3 ( TID3 ) ,.TID2 ( TID2 )
     ,.TID1 ( TID1 ) ,.TID0 ( TID0 ) ,.TESINST ( TESINST ) ,.BBTESINST ( BBTESINST )
     ,.PTESINST ( PTESINST ) ,.OPTFLMEM ( OPTFLMEM ) ,.OPTMDUMP ( OPTMDUMP )
     ,.SPRGMOD ( SPRGMOD ) ,.TESTMOD ( TESTMOD ) ,.TMODDFT ( TESTMOD )
     ,.READ ( READ ) ,.TESDBT ( TESDBT ) ,.SCANMODE ( SCANMODE ) ,.SELRO1 ( SELRO1 )
     ,.TA17 ( TA17 ) ,.TA16 ( TA16 ) ,.TA15 ( TA15 ) ,.TA14 ( TA14 ) ,.TA13 ( TA13 )
     ,.TA12 ( TA12 ) ,.TA11 ( TA11 ) ,.TA10 ( TA10 ) ,.TA9 ( TA9 ) ,.TA8 ( TA8 )
     ,.TA7 ( TA7 ) ,.TA6 ( TA6 ) ,.TA5 ( TA5 ) ,.TA4 ( TA4 ) ,.TA2 ( TA2 )
     ,.TA1 ( TA1 ) ,.TA0 ( TA0 ) ,.FRQSEL4 ( FRQSEL4 ) ,.FRQSEL3 ( FRQSEL3 )
     ,.FRQSEL2 ( FRQSEL2 ) ,.FRQSEL1 ( FRQSEL1 ) ,.FRQSEL0 ( FRQSEL0 )
     ,.RLOWSPY ( RLOWSPY ) ,.LOWPOWER ( LOWPOWER ) ,.MODEFNOP ( MODEFNOP )
     ,.TPIDSEL ( TPIDSEL ) ,.CTRIM6 ( CTRIM6 ) ,.CTRIM5 ( CTRIM5 ) ,.CTRIM4 ( CTRIM4 )
     ,.CTRIM3 ( CTRIM3 ) ,.CTRIM2 ( CTRIM2 ) ,.CTRIM1 ( CTRIM1 ) ,.CTRIM0 ( CTRIM0 )
     ,.WTRIM2 ( WTRIM2 ) ,.WTRIM1 ( WTRIM1 ) ,.WTRIM0 ( WTRIM0 ) ,.FTRIM5 ( FTRIM5 )
     ,.FTRIM4 ( FTRIM4 ) ,.FTRIM3 ( FTRIM3 ) ,.FTRIM2 ( FTRIM2 ) ,.FTRIM1 ( FTRIM1 )
     ,.FTRIM0 ( FTRIM0 ) ,.RTRIM5 ( RTRIM5 ) ,.RTRIM4 ( RTRIM4 ) ,.RTRIM3 ( RTRIM3 )
     ,.RTRIM2 ( RTRIM2 ) ,.RTRIM1 ( RTRIM1 ) ,.RTRIM0 ( RTRIM0 ) ,.BGRT10 ( BGRT10 )
     ,.BGRT9 ( BGRT9 ) ,.BGRT8 ( BGRT8 ) ,.BGRT7 ( BGRT7 ) ,.BGRT6 ( BGRT6 )
     ,.BGRT5 ( BGRT5 ) ,.BGRT4 ( BGRT4 ) ,.BGRT3 ( BGRT3 ) ,.BGRT2 ( BGRT2 )
     ,.BGRT1 ( BGRT1 ) ,.BGRT0 ( BGRT0 ) ,.OPBOEN ( OPBOEN ) ,.BBNVM1 ( BBNVM1 )
     ,.BBNVM2 ( BBNVM2 ) ,.PSEL4 ( PSELCIB4 ) ,.CSPDTFLG ( CSPDTFLP ) ,.CKSMER ( CKSMER )
     ,.CFNSD9 ( CFNSD9 ) ,.CFNSD8 ( CFNSD8 ) ,.CFNSD7 ( CFNSD7 ) ,.CFNSD6 ( CFNSD6 )
     ,.CFNSD5 ( CFNSD5 ) ,.CFNSD4 ( CFNSD4 ) ,.CFNSD3 ( CFNSD3 ) ,.CFNSD2 ( CFNSD2 )
     ,.CFNSD1 ( CFNSD1 ) ,.CFNSD0 ( CFNSD0 ) ,.WWR ( WWR ) ,.FSWE9 ( FSWE9 )
     ,.FSWE8 ( FSWE8 ) ,.FSWE7 ( FSWE7 ) ,.FSWE6 ( FSWE6 ) ,.FSWE5 ( FSWE5 )
     ,.FSWE4 ( FSWE4 ) ,.FSWE3 ( FSWE3 ) ,.FSWE2 ( FSWE2 ) ,.FSWE1 ( FSWE1 )
     ,.FSWE0 ( FSWE0 ) ,.CIBRESRQ ( CIBRESRQ ) ,.SELTAF ( SELTAF ) ,.CECCE ( CECCE )
     ,.TMSPMD ( ICETMSPMD ) ,.BTFLG ( BTFLG ) ,.TRMRD1CK ( TRMRD1CK ) ,.TRMRD2CK ( TRMRD2CK )
     ,.BRSAM ( BRSAM ) ,.FSPR ( FSPR ) ,.RDPR ( RDPR ) ,.WRPR ( WRPR )
     ,.SEPR ( SEPR ) ,.BTPR ( BTPR ) ,.BTBLS1 ( BTBLS1 ) ,.BTBLS0 ( BTBLS0 )
     ,.FPSER2 ( FPSER2 ) ,.FPSER1 ( FPSER1 ) ,.FPSER0 ( FPSER0 ) ,.FPWWR2 ( FPWWR2 )
     ,.FPWWR1 ( FPWWR1 ) ,.FPWWR0 ( FPWWR0 ) ,.FPERTY7 ( FPERTY7 ) ,.FPERTY6 ( FPERTY6 )
     ,.FPERTY5 ( FPERTY5 ) ,.FPERTY4 ( FPERTY4 ) ,.FPERTY3 ( FPERTY3 )
     ,.FPERTY2 ( FPERTY2 ) ,.FPERTY1 ( FPERTY1 ) ,.FPERTY0 ( FPERTY0 )
     ,.FPWRTY7 ( FPWRTY7 ) ,.FPWRTY6 ( FPWRTY6 ) ,.FPWRTY5 ( FPWRTY5 )
     ,.FPWRTY4 ( FPWRTY4 ) ,.FPWRTY3 ( FPWRTY3 ) ,.FPWRTY2 ( FPWRTY2 )
     ,.FPWRTY1 ( FPWRTY1 ) ,.FPWRTY0 ( FPWRTY0 ) ,.FPECC3 ( FPECC3 ) ,.FPECC2 ( FPECC2 )
     ,.FPECC1 ( FPECC1 ) ,.FPECC0 ( FPECC0 ) ,.R0FLAGZ ( R0FLAGZ ) ,.R1FLAGZ ( R1FLAGZ )
     ,.R0A7 ( R0A7 ) ,.R1A3 ( R1A3 ) ,.R0A6 ( R0A6 ) ,.R1A2 ( R1A2 ) ,.R0A5 ( R0A5 )
     ,.R1A1 ( R1A1 ) ,.R0A4 ( R0A4 ) ,.R1A0 ( R1A0 ) ,.R0A3 ( R0A3 ) ,.R0A2 ( R0A2 )
     ,.R0A1 ( R0A1 ) ,.R0A0 ( R0A0 ) ,.R1A7 ( R1A7 ) ,.R1A6 ( R1A6 ) ,.R1A5 ( R1A5 )
     ,.R1A4 ( R1A4 ) ,.ICENOECC ( ICENOECC ) ,.SLECCOFF ( SLECCOFF ) ,.ECCER ( ECCER )
     ,.FMULTIEN ( FMULTIEN ) ,.OSCNOSTP ( OSCNOSTP ) ,.POSCNOST ( POSCNOST )
     ,.POSCOUTE ( POSCOUTE ) ,.CPT ( CPT ) ,.TESTRMRD ( TESTRMRD ) ,.HIOMSK ( HIOMSK )
     ,.SCANCLK ( SCANCLK ) ,.TFLSTOPC ( TFLSTOPC ) ,.AisRSEQ ( AisRSEQ )
     ,.RDSETUP ( RDSETUP ) ,.FLROACT ( FLROACT ) ,.FRQ4EN ( FRQ4EN ) ,.PSYSRESB ( PSYSRESB )
     ,.CHMOD ( CHMOD ) ,.GOFIRMR ( GOFIRMR )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_soft/qlk0rcibdm3sf1v1_mf3_1.20/_library/101015/qlk0rcibdm3sf1v1.hdl
  QLK0RCIBDM3SF1V1 cibd (
    .PENABLE ( PENABLE ) ,.PWRITE ( PWRITE ) ,.PSEL1 ( PSELCIBD ) ,.PADDR1 ( PADDR1 )
     ,.PWDATA7 ( MDW7 ) ,.PWDATA4 ( MDW4 ) ,.PWDATA3 ( MDW3 ) ,.PWDATA0 ( MDW0 )
     ,.PRDATA15 ( PRDCID15 ) ,.PRDATA14 ( PRDCID14 ) ,.PRDATA13 ( PRDCID13 )
     ,.PRDATA12 ( PRDCID12 ) ,.PRDATA11 ( PRDCID11 ) ,.PRDATA10 ( PRDCID10 )
     ,.PRDATA9 ( PRDCID9 ) ,.PRDATA8 ( PRDCID8 ) ,.SELTADF ( SELTADF )
     ,.PRDATA7 ( PRDCID7 ) ,.PRDATA6 ( PRDCID6 ) ,.PRDATA5 ( PRDCID5 )
     ,.PRDATA4 ( PRDCID4 ) ,.PRDATA3 ( PRDCID3 ) ,.PRDATA2 ( PRDCID2 )
     ,.PRDATA1 ( PRDCID1 ) ,.PRDATA0 ( PRDCID0 ) ,.BASECKHS ( BASECKHS )
     ,.RESETB ( RESETB ) ,.SCANCLK ( SCANCLK ) ,.RESB ( RESB ) ,.MA13 ( MA13 )
     ,.MA12 ( MA12 ) ,.MA11 ( MA11 ) ,.MA10 ( MA10 ) ,.MA9 ( MA9 ) ,.MA8 ( MA8 )
     ,.MA7 ( MA7 ) ,.MA6 ( MA6 ) ,.MA5 ( MA5 ) ,.MA4 ( MA4 ) ,.MA3 ( MA3 )
     ,.MA2 ( MA2 ) ,.MA1 ( MA1 ) ,.MA0 ( MA0 ) ,.MDR15 ( MDRCID15 ) ,.MDR14 ( MDRCID14 )
     ,.MDR13 ( MDRCID13 ) ,.MDR12 ( MDRCID12 ) ,.MDR11 ( MDRCID11 ) ,.MDR10 ( MDRCID10 )
     ,.MDR9 ( MDRCID9 ) ,.MDR8 ( MDRCID8 ) ,.MDR7 ( MDRCID7 ) ,.MDR6 ( MDRCID6 )
     ,.MDR5 ( MDRCID5 ) ,.MDR4 ( MDRCID4 ) ,.MDR3 ( MDRCID3 ) ,.MDR2 ( MDRCID2 )
     ,.MDR1 ( MDRCID1 ) ,.MDR0 ( MDRCID0 ) ,.SLDFLASH ( SLDFLASH ) ,.FHLTST ( FHLTST )
     ,.FSTPST ( FSTPST ) ,.SUB ( SUB ) ,.AF13 ( AF13 ) ,.AF12 ( AF12 )
     ,.AF11 ( AF11 ) ,.AF10 ( AF10 ) ,.AF9 ( AF9 ) ,.DA7 ( DA7 ) ,.AF8 ( AF8 )
     ,.DA6 ( DA6 ) ,.AF7 ( AF7 ) ,.DA5 ( DA5 ) ,.AF6 ( AF6 ) ,.DA4 ( DA4 )
     ,.AF5 ( AF5 ) ,.DA3 ( DA3 ) ,.AF4 ( AF4 ) ,.DA2 ( DA2 ) ,.AF3 ( AF3 )
     ,.DA1 ( DA1 ) ,.AF2 ( AF2 ) ,.DA0 ( DA0 ) ,.AF1 ( AF1 ) ,.AF0 ( AF0 )
     ,.DFLRO11 ( DFLRO11 ) ,.DFLRO10 ( DFLRO10 ) ,.DFLRO9 ( DFLRO9 ) ,.DFLRO8 ( DFLRO8 )
     ,.DFLRO7 ( DFLRO7 ) ,.DFLRO6 ( DFLRO6 ) ,.DFLRO5 ( DFLRO5 ) ,.DFLRO4 ( DFLRO4 )
     ,.DFLRO3 ( DFLRO3 ) ,.DFLRO2 ( DFLRO2 ) ,.DFLRO1 ( DFLRO1 ) ,.DFLRO0 ( DFLRO0 )
     ,.SACEEN ( SACEEN ) ,.DCE0 ( DCE0 ) ,.DA13 ( DA13 ) ,.DA12 ( DA12 )
     ,.DA11 ( DA11 ) ,.DA10 ( DA10 ) ,.DA9 ( DA9 ) ,.DA8 ( DA8 ) ,.DRO011 ( DRO011 )
     ,.DRO010 ( DRO010 ) ,.DRO09 ( DRO09 ) ,.DRO08 ( DRO08 ) ,.DRO07 ( DRO07 )
     ,.DRO06 ( DRO06 ) ,.DRO05 ( DRO05 ) ,.DRO04 ( DRO04 ) ,.DRO03 ( DRO03 )
     ,.DRO02 ( DRO02 ) ,.DRO01 ( DRO01 ) ,.DRO00 ( DRO00 ) ,.DCLKSEL1 ( DCLKSEL1 )
     ,.DSRCUT ( DSRCUT ) ,.DFLSTOP ( DFLSTOP ) ,.OPTMDUMP ( OPTMDUMP )
     ,.TESTMOD ( TESTMOD ) ,.TMODDFT ( TESTMOD ) ,.TESDBT ( TESDBT ) ,.SCANMODE ( SCANMODE )
     ,.TA13 ( TA13 ) ,.TA12 ( TA12 ) ,.TA11 ( TA11 ) ,.TA10 ( TA10 ) ,.TA9 ( TA9 )
     ,.TA8 ( TA8 ) ,.TA7 ( TA7 ) ,.TA6 ( TA6 ) ,.TA5 ( TA5 ) ,.TA4 ( TA4 )
     ,.TA3 ( TA3 ) ,.TA2 ( TA2 ) ,.TA1 ( TA1 ) ,.TA0 ( TA0 ) ,.DECCE ( DECCE )
     ,.EEEMD ( EEEMD ) ,.DFLEN ( DFLEN ) ,.DRDCLK ( DRDCLK ) ,.DRDCLKC1 ( DRDCLKC1 )
     ,.ICENOECC ( ICENOECC ) ,.OPTDFL ( OPTDFL ) ,.SLECCOFF ( SLECCOFF )
     ,.DECCER ( DECCER ) ,.STDWAIT ( STDWAIT ) ,.TFLSTOPD ( TFLSTOPD )
     ,.AisRSEQ ( AisRSEQ ) ,.RDSETUP ( RDSETUP ) ,.BASECK ( BASECK )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_soft/qlk0rfcbm3sf1v1_rtl_v1.20_LR2.0.01_20100823/_misc/QLK0RFCBM3SF1V1.v
  QLK0RFCBM3SF1V1 fcb (
    .TESTMOD ( TESTMOD ) ,.BTBLS1 ( BTBLS1 ) ,.BTBLS0 ( BTBLS0 ) ,.FSWE9 ( FSWE9 )
     ,.FSWE8 ( FSWE8 ) ,.FSWE7 ( FSWE7 ) ,.FSWE6 ( FSWE6 ) ,.IREFT ( IREFT )
     ,.FSWE5 ( FSWE5 ) ,.FSWE4 ( FSWE4 ) ,.FSWE3 ( FSWE3 ) ,.FSWE2 ( FSWE2 )
     ,.MRG12 ( MRG12 ) ,.FSWE1 ( FSWE1 ) ,.MRG11 ( MRG11 ) ,.FSWE0 ( FSWE0 )
     ,.MRG10 ( MRG10 ) ,.FSWS9 ( FSWS9 ) ,.FSWS8 ( FSWS8 ) ,.FSWS7 ( FSWS7 )
     ,.FSWS6 ( FSWS6 ) ,.FSWS5 ( FSWS5 ) ,.FSWS4 ( FSWS4 ) ,.FSWS3 ( FSWS3 )
     ,.FSWS2 ( FSWS2 ) ,.FSWEN ( FSWEN ) ,.FSWS1 ( FSWS1 ) ,.FSWS0 ( FSWS0 )
     ,.FLSPM ( FLSPM ) ,.EEEMD ( EEEMD ) ,.LOWSPY ( LOWSPY ) ,.CWEE ( CWEE )
     ,.SCANMODE ( SCANMODE ) ,.EXCHEN ( EXCHEN ) ,.SECEN ( SECEN ) ,.FPSER2 ( FPSER2 )
     ,.FPSER1 ( FPSER1 ) ,.FPSER0 ( FPSER0 ) ,.FPWWR2 ( FPWWR2 ) ,.FPWWR1 ( FPWWR1 )
     ,.FPWWR0 ( FPWWR0 ) ,.FPWRTY7 ( FPWRTY7 ) ,.FPWRTY6 ( FPWRTY6 ) ,.FPWRTY5 ( FPWRTY5 )
     ,.FPWRTY4 ( FPWRTY4 ) ,.FPWRTY3 ( FPWRTY3 ) ,.FPWRTY2 ( FPWRTY2 )
     ,.FPWRTY1 ( FPWRTY1 ) ,.FPWRTY0 ( FPWRTY0 ) ,.FPERTY7 ( FPERTY7 )
     ,.FPERTY6 ( FPERTY6 ) ,.FPERTY5 ( FPERTY5 ) ,.FPERTY4 ( FPERTY4 )
     ,.FPERTY3 ( FPERTY3 ) ,.FPERTY2 ( FPERTY2 ) ,.FPERTY1 ( FPERTY1 )
     ,.FPERTY0 ( FPERTY0 ) ,.FPECC3 ( FPECC3 ) ,.FPECC2 ( FPECC2 ) ,.FPECC1 ( FPECC1 )
     ,.FPECC0 ( FPECC0 ) ,.CECCE ( CECCE ) ,.DECCE ( DECCE ) ,.INTFL ( INTFL )
     ,.STDWAIT ( STDWAIT ) ,.TMBTSEL ( TMBTSEL ) ,.TMSPMD ( TMSPMD ) ,.EXCH ( EXCH )
     ,.FSPR ( FSPR ) ,.RDPR ( RDPR ) ,.WRPR ( WRPR ) ,.CEPR ( CEPR ) ,.SEPR ( SEPR )
     ,.BTPR ( BTPR ) ,.BTFLG ( BTFLG ) ,.DDIS ( DDIS ) ,.DW33 ( DW33 )
     ,.DW25 ( DW25 ) ,.DW17 ( DW17 ) ,.DREAD ( DREAD ) ,.DMRG00 ( DMRG00 )
     ,.DMRG01 ( DMRG01 ) ,.DMRG10 ( DMRG10 ) ,.DMRG11 ( DMRG11 ) ,.DMRG12 ( DMRG12 )
     ,.DSER ( DSER ) ,.DWWR ( DWWR ) ,.DCER ( DCER ) ,.PSEL2 ( PSELFCB2 )
     ,.PSEL1 ( PSELFCB1 ) ,.PADDR4 ( PADDR4 ) ,.PADDR3 ( PADDR3 ) ,.PADDR2 ( PADDR2 )
     ,.PADDR1 ( PADDR1 ) ,.PADDR0 ( PADDR0 ) ,.PWDATA15 ( MDW15 ) ,.PWDATA14 ( MDW14 )
     ,.PWDATA13 ( MDW13 ) ,.PWDATA12 ( MDW12 ) ,.PWDATA11 ( MDW11 ) ,.PWDATA10 ( MDW10 )
     ,.PWDATA9 ( MDW9 ) ,.PWDATA8 ( MDW8 ) ,.PWDATA7 ( MDW7 ) ,.PWDATA6 ( MDW6 )
     ,.PWDATA5 ( MDW5 ) ,.PWDATA4 ( MDW4 ) ,.PWDATA3 ( MDW3 ) ,.PWDATA2 ( MDW2 )
     ,.PWDATA1 ( MDW1 ) ,.PWDATA0 ( MDW0 ) ,.PRDATA15 ( PRDFCB15 ) ,.PRDATA14 ( PRDFCB14 )
     ,.PRDATA13 ( PRDFCB13 ) ,.PRDATA12 ( PRDFCB12 ) ,.PRDATA11 ( PRDFCB11 )
     ,.PRDATA10 ( PRDFCB10 ) ,.PRDATA9 ( PRDFCB9 ) ,.PRDATA8 ( PRDFCB8 )
     ,.PRDATA7 ( PRDFCB7 ) ,.PRDATA6 ( PRDFCB6 ) ,.PRDATA5 ( PRDFCB5 )
     ,.PRDATA4 ( PRDFCB4 ) ,.PRDATA3 ( PRDFCB3 ) ,.PRDATA2 ( PRDFCB2 )
     ,.PRDATA1 ( PRDFCB1 ) ,.PRDATA0 ( PRDFCB0 ) ,.PWRITE ( PWRITE ) ,.PRESETZ ( RESETB )
     ,.PENABLE ( PENABLE ) ,.FLMEMTES ( FLMEMTES ) ,.DIS ( DIS ) ,.DW7 ( DW7 )
     ,.READ ( READ ) ,.MRG00 ( MRG00 ) ,.MRG01 ( MRG01 ) ,.WWR ( WWR )
     ,.MSWR ( MSWR ) ,.CER ( CER ) ,.SER ( SER ) ,.EXER ( EXER ) ,.STCHK ( STCHK )
     ,.IONCHK1 ( IONCHK1 ) ,.RDT ( RDT ) ,.RDMRG1 ( RDMRG1 ) ,.RDMRG0 ( RDMRG0 )
     ,.RDMRGC ( RDMRGC ) ,.WDT1 ( WDT1 ) ,.WDT2 ( WDT2 ) ,.WDT3 ( WDT3 )
     ,.WDT4 ( WDT4 ) ,.CPBT ( CPBT ) ,.SACEEN ( SACEEN ) ,.CPT ( CPT )
     ,.EXTVPP2 ( EXTVPP2 ) ,.EXTVPP1 ( EXTVPP1 ) ,.MEOC ( MEOC ) ,.MEOR ( MEOR )
     ,.BEU2 ( BEU2 ) ,.BEU1 ( BEU1 ) ,.BEU0 ( BEU0 ) ,.MODIDIS ( MODIDIS )
     ,.TFWEPR ( pull_up48 ) ,.MUTEST ( MUTEST ) ,.EXA ( PEXA ) ,.WED ( WED )
     ,.DWED ( DWED ) ,.ONBD ( SPRGMOD ) ,.DFLRO11 ( DFLRO11 ) ,.DFLRO10 ( DFLRO10 )
     ,.DFLRO9 ( DFLRO9 ) ,.DFLRO8 ( DFLRO8 ) ,.DFLRO7 ( DFLRO7 ) ,.DFLRO6 ( DFLRO6 )
     ,.DFLRO5 ( DFLRO5 ) ,.DFLRO4 ( DFLRO4 ) ,.DFLRO3 ( DFLRO3 ) ,.DFLRO2 ( DFLRO2 )
     ,.DFLRO1 ( DFLRO1 ) ,.DFLRO0 ( DFLRO0 ) ,.FLRO37 ( FLRO37 ) ,.FLRO29 ( FLRO29 )
     ,.FLRO36 ( FLRO36 ) ,.FLRO28 ( FLRO28 ) ,.FLRO35 ( FLRO35 ) ,.FLRO27 ( FLRO27 )
     ,.FLRO19 ( FLRO19 ) ,.FLRO34 ( FLRO34 ) ,.FLRO26 ( FLRO26 ) ,.FLRO18 ( FLRO18 )
     ,.FLRO33 ( FLRO33 ) ,.FLRO25 ( FLRO25 ) ,.FLRO17 ( FLRO17 ) ,.FLRO32 ( FLRO32 )
     ,.FLRO24 ( FLRO24 ) ,.FLRO16 ( FLRO16 ) ,.FLRO31 ( FLRO31 ) ,.FLRO23 ( FLRO23 )
     ,.FLRO15 ( FLRO15 ) ,.FLRO30 ( FLRO30 ) ,.FLRO22 ( FLRO22 ) ,.FLRO14 ( FLRO14 )
     ,.FLRO21 ( FLRO21 ) ,.FLRO13 ( FLRO13 ) ,.FLRO20 ( FLRO20 ) ,.FLRO12 ( FLRO12 )
     ,.FLRO11 ( FLRO11 ) ,.FLRO10 ( FLRO10 ) ,.FLRO9 ( FLRO9 ) ,.FLRO8 ( FLRO8 )
     ,.FLRO7 ( FLRO7 ) ,.FLRO6 ( FLRO6 ) ,.FLRO5 ( FLRO5 ) ,.FLRO4 ( FLRO4 )
     ,.FLRO3 ( FLRO3 ) ,.FLRO2 ( FLRO2 ) ,.FLRO1 ( FLRO1 ) ,.FLRO0 ( FLRO0 )
     ,.DW37 ( DW37 ) ,.DW29 ( DW29 ) ,.DW36 ( DW36 ) ,.DW28 ( DW28 ) ,.DW35 ( DW35 )
     ,.DW27 ( DW27 ) ,.DW19 ( DW19 ) ,.DW34 ( DW34 ) ,.DW26 ( DW26 ) ,.DW18 ( DW18 )
     ,.DW32 ( DW32 ) ,.DW24 ( DW24 ) ,.DW16 ( DW16 ) ,.DW31 ( DW31 ) ,.DW23 ( DW23 )
     ,.DW15 ( DW15 ) ,.DW30 ( DW30 ) ,.DW22 ( DW22 ) ,.DW14 ( DW14 ) ,.DW21 ( DW21 )
     ,.DW13 ( DW13 ) ,.DW20 ( DW20 ) ,.DW12 ( DW12 ) ,.DW11 ( DW11 ) ,.DW10 ( DW10 )
     ,.DW9 ( DW9 ) ,.DW8 ( DW8 ) ,.DW6 ( DW6 ) ,.DW5 ( DW5 ) ,.DW4 ( DW4 )
     ,.DW3 ( DW3 ) ,.DW2 ( DW2 ) ,.DW1 ( DW1 ) ,.DW0 ( DW0 ) ,.FCLK1 ( FCLK1 )
     ,.FCLK2 ( FCLK2 ) ,.RDCLKP1 ( RDCLKP1 ) ,.PROGI ( PROGI ) ,.AF19 ( AF19 )
     ,.AF18 ( AF18 ) ,.AF17 ( AF17 ) ,.AF16 ( AF16 ) ,.AF15 ( AF15 ) ,.AF14 ( AF14 )
     ,.AF13 ( AF13 ) ,.AF12 ( AF12 ) ,.AF11 ( AF11 ) ,.AF10 ( AF10 ) ,.AF9 ( AF9 )
     ,.AF8 ( AF8 ) ,.AF7 ( AF7 ) ,.AF6 ( AF6 ) ,.AF5 ( AF5 ) ,.AF4 ( AF4 )
     ,.AF3 ( AF3 ) ,.AF2 ( AF2 ) ,.AF1 ( AF1 ) ,.AF0 ( AF0 ) ,.SSEQBRK ( SVSTOP )
     ,.ICENOECC ( ICENOECC ) ,.ICEFLERR ( ICEFLERR ) ,.PCLK ( PCLKFCB )
     ,.VCEQ ( VCEQ )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/qlk0rwwdt1v2_v2.20_LR3.0.01_20100820/_library/QLK0RWWDT1V2.v
  QLK0RWWDT1V2 wwdt (
    .PCLKRW ( PCLKRW ) ,.PRESETZ ( PRESWDTZ ) ,.PWDATA15 ( MDW15 ) ,.PWDATA14 ( MDW14 )
     ,.PWDATA13 ( MDW13 ) ,.PWDATA12 ( MDW12 ) ,.PWDATA11 ( MDW11 ) ,.PWDATA10 ( MDW10 )
     ,.PWDATA9 ( MDW9 ) ,.OPWDCS1 ( OPWDCS1 ) ,.PWDATA8 ( MDW8 ) ,.OPWDCS0 ( OPWDCS0 )
     ,.PRDATA15 ( PRDWDT15 ) ,.PRDATA12 ( PRDWDT12 ) ,.PRDATA11 ( PRDWDT11 )
     ,.PRDATA9 ( PRDWDT9 ) ,.PWRITE ( PWRITE ) ,.PENABLE ( PENABLE ) ,.PSEL ( PSELWWDT )
     ,.WDEN ( WDEN ) ,.OPWDCS2 ( OPWDCS2 ) ,.OPWDWS1 ( OPWDWS1 ) ,.OPWDWS0 ( OPWDWS0 )
     ,.OPWDINT ( OPWDINT ) ,.OPWDSTBY ( OPWDSTBY ) ,.CPUSTART ( CPUSTART )
     ,.SCANMODE ( SCANMODE ) ,.SVMOD ( SVSTOP ) ,.SPRGMOD ( SPRGMOD ) ,.WDTRES ( WDTRES )
     ,.INTWWDT ( INTWWDT ) ,.WDTCLK ( R15KOUT ) ,.WDTTESCK ( WDTTESCK )
     ,.WDTTEN ( OPTBCT ) ,.WDTMON ( WDTMON )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/qlk0rrtc0v3_v3.10_LR3.0.04_20100721/_library/QLK0RRTC0V3.v
  QLK0RRTC0V3 rtc (
    .SCANMODE ( SCANMODE ) ,.RT0LPM ( RT0LPM ) ,.PCLK ( PCLKRTC ) ,.RTCRESB ( PRESRTCZ )
     ,.PRESETZ ( PRESRTCZ ) ,.RTCCLK ( RTCCLK ) ,.INTRCLK ( INTRCLK ) ,.CKSEL ( CKSEL )
     ,.RT0TEN ( OPTBCT ) ,.SVMOD ( SVPERI0 ) ,.PADDR3 ( PADDR3 ) ,.PADDR2 ( PADDR2 )
     ,.PADDR1 ( PADDR1 ) ,.PADDR0 ( PADDR0 ) ,.PWDATA15 ( MDW15 ) ,.PWDATA14 ( MDW14 )
     ,.PWDATA13 ( MDW13 ) ,.PWDATA12 ( MDW12 ) ,.PWDATA11 ( MDW11 ) ,.PWDATA10 ( MDW10 )
     ,.PWDATA9 ( MDW9 ) ,.PWDATA8 ( MDW8 ) ,.PWDATA7 ( MDW7 ) ,.PWDATA6 ( MDW6 )
     ,.PWDATA5 ( MDW5 ) ,.PWDATA4 ( MDW4 ) ,.PWDATA3 ( MDW3 ) ,.PWDATA2 ( MDW2 )
     ,.PWDATA1 ( MDW1 ) ,.PWDATA0 ( MDW0 ) ,.PRDATA15 ( PRDRTC15 ) ,.PRDATA14 ( PRDRTC14 )
     ,.PRDATA13 ( PRDRTC13 ) ,.PRDATA12 ( PRDRTC12 ) ,.PRDATA11 ( PRDRTC11 )
     ,.PRDATA10 ( PRDRTC10 ) ,.PRDATA9 ( PRDRTC9 ) ,.PRDATA8 ( PRDRTC8 )
     ,.PRDATA7 ( PRDRTC7 ) ,.PRDATA6 ( PRDRTC6 ) ,.PRDATA5 ( PRDRTC5 )
     ,.PRDATA4 ( PRDRTC4 ) ,.PRDATA3 ( PRDRTC3 ) ,.PRDATA2 ( PRDRTC2 )
     ,.PRDATA1 ( PRDRTC1 ) ,.PRDATA0 ( PRDRTC0 ) ,.PWRITE ( PWRITE ) ,.PENABLE ( PENABLE )
     ,.PSEL ( PSELRTC ) ,.INTRTC ( INTRTC ) ,.INTRTCI ( INTRTCI ) ,.CLK1HZ ( CLK1HZ )
     ,.RT0MON0 ( RT0MON0 ) ,.RT0MON1 ( RT0MON1 )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_soft/qlk0rcrc0v1_mf3_v1.00/_library/100412/qlk0rcrc0v1.hdl
  QLK0RCRC0V1 crc (
    .PWRITE ( PWRITE ) ,.PSELCRC ( PSELCRC ) ,.PENABLE ( PENABLE ) ,.PWDATA15 ( MDW15 )
     ,.PWDATA14 ( MDW14 ) ,.PWDATA13 ( MDW13 ) ,.PWDATA12 ( MDW12 ) ,.PWDATA11 ( MDW11 )
     ,.PWDATA10 ( MDW10 ) ,.PWDATA9 ( MDW9 ) ,.PWDATA8 ( MDW8 ) ,.PWDATA7 ( MDW7 )
     ,.PWDATA6 ( MDW6 ) ,.PWDATA5 ( MDW5 ) ,.PWDATA4 ( MDW4 ) ,.PWDATA3 ( MDW3 )
     ,.PWDATA2 ( MDW2 ) ,.PWDATA1 ( MDW1 ) ,.PWDATA0 ( MDW0 ) ,.PRDATA15 ( PRDCRC15 )
     ,.PRDATA14 ( PRDCRC14 ) ,.PRDATA13 ( PRDCRC13 ) ,.PRDATA12 ( PRDCRC12 )
     ,.PRDATA11 ( PRDCRC11 ) ,.PRDATA10 ( PRDCRC10 ) ,.PRDATA9 ( PRDCRC9 )
     ,.PRDATA8 ( PRDCRC8 ) ,.PRDATA7 ( PRDCRC7 ) ,.PRDATA6 ( PRDCRC6 )
     ,.PRDATA5 ( PRDCRC5 ) ,.PRDATA4 ( PRDCRC4 ) ,.PRDATA3 ( PRDCRC3 )
     ,.PRDATA2 ( PRDCRC2 ) ,.PRDATA1 ( PRDCRC1 ) ,.PRDATA0 ( PRDCRC0 )
     ,.PADDR1 ( PADDR1 ) ,.PADDR0 ( PADDR0 ) ,.BASECK ( BASECKHS ) ,.RESB ( RESB )
     ,.PCLKRW ( PCLKRW )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/_ice/_macro/_sss/maw/100910/qlk0rmaw0v1.hdl
  QLK0RMAW0V1 maw0 (
    .PENABLE ( PENABLE ) ,.PWRITE ( PWRITE ) ,.PSEL ( PSELMAW ) ,.PADDR2 ( PADDR2 )
     ,.PADDR1 ( PADDR1 ) ,.PADDR0 ( PADDR0 ) ,.PWDATA15 ( MDW15 ) ,.PWDATA14 ( MDW14 )
     ,.PWDATA13 ( MDW13 ) ,.PWDATA12 ( MDW12 ) ,.PWDATA11 ( MDW11 ) ,.PWDATA10 ( MDW10 )
     ,.PWDATA9 ( MDW9 ) ,.PWDATA8 ( MDW8 ) ,.PWDATA7 ( MDW7 ) ,.BASECK ( BASECK )
     ,.RESB ( RESB ) ,.SYSRESB ( SYSRESB ) ,.PC19 ( MONPC19 ) ,.PC18 ( MONPC18 )
     ,.PC17 ( MONPC17 ) ,.PC16 ( MONPC16 ) ,.PC15 ( MONPC15 ) ,.PC14 ( MONPC14 )
     ,.PC13 ( MONPC13 ) ,.PC12 ( MONPC12 ) ,.PC11 ( MONPC11 ) ,.PA19 ( PA19 )
     ,.PC10 ( MONPC10 ) ,.PA18 ( PA18 ) ,.PC9 ( MONPC9 ) ,.PC8 ( MONPC8 )
     ,.PC7 ( MONPC7 ) ,.PC6 ( MONPC6 ) ,.PC5 ( MONPC5 ) ,.PA9 ( PA9 ) ,.PC4 ( MONPC4 )
     ,.PA8 ( PA8 ) ,.PC3 ( MONPC3 ) ,.PA7 ( PA7 ) ,.PC2 ( MONPC2 ) ,.PA6 ( PA6 )
     ,.PC1 ( MONPC1 ) ,.PA5 ( PA5 ) ,.PC0 ( MONPC0 ) ,.PA4 ( PA4 ) ,.PA17 ( PA17 )
     ,.PA16 ( PA16 ) ,.PA15 ( PA15 ) ,.PA14 ( PA14 ) ,.PA13 ( PA13 ) ,.PA12 ( PA12 )
     ,.PA11 ( PA11 ) ,.PA10 ( PA10 ) ,.PA3 ( PA3 ) ,.PA2 ( PA2 ) ,.MA15 ( MONMA15 )
     ,.MA14 ( MONMA14 ) ,.MA13 ( MONMA13 ) ,.MA12 ( MONMA12 ) ,.MA11 ( MONMA11 )
     ,.MA10 ( MONMA10 ) ,.MA9 ( MONMA9 ) ,.MA8 ( MONMA8 ) ,.MA7 ( MONMA7 )
     ,.MA6 ( MONMA6 ) ,.MA5 ( MONMA5 ) ,.MA4 ( MONMA4 ) ,.MA3 ( MONMA3 )
     ,.MA2 ( MONMA2 ) ,.MA1 ( MONMA1 ) ,.MA0 ( MONMA0 ) ,.CPURD ( CPURD )
     ,.CPUWR ( CPUWR ) ,.SLFLASH ( SLFLASH ) ,.SLMEM ( SLMEM ) ,.FLREAD ( FLREAD )
     ,.FCHRAM ( FCHRAM ) ,.FLSIZE3 ( FLSIZE3 ) ,.FLSIZE2 ( FLSIZE2 ) ,.FLSIZE1 ( FLSIZE1 )
     ,.FLSIZE0 ( FLSIZE0 ) ,.RAMSIZE7 ( pull_up51 ) ,.RAMSIZE6 ( pull_up52 )
     ,.RAMSIZE5 ( pull_up53 ) ,.RAMSIZE4 ( pull_down12 ) ,.RAMSIZE3 ( pull_up54 )
     ,.RAMSIZE2 ( pull_up55 ) ,.RAMSIZE1 ( pull_up56 ) ,.RAMSIZE0 ( pull_up57 )
     ,.BFSIZE3 ( BFSIZE3 ) ,.BFSIZE2 ( BFSIZE2 ) ,.BFSIZE1 ( BFSIZE1 )
     ,.BFSIZE0 ( BFSIZE0 ) ,.BMSIZE3 ( BMSIZE3 ) ,.BMSIZE2 ( BMSIZE2 )
     ,.BMSIZE1 ( BMSIZE1 ) ,.BMSIZE0 ( BMSIZE0 ) ,.DMARD ( DMARD ) ,.DMAWR ( DMAWR )
     ,.PBFA ( pull_up50 ) ,.CFNSD9 ( CFNSD9 ) ,.CFNSD8 ( CFNSD8 ) ,.CFNSD7 ( CFNSD7 )
     ,.CFNSD6 ( CFNSD6 ) ,.CFNSD5 ( CFNSD5 ) ,.CFNSD4 ( CFNSD4 ) ,.CFNSD3 ( CFNSD3 )
     ,.CFNSD2 ( CFNSD2 ) ,.CFNSD1 ( CFNSD1 ) ,.CFNSD0 ( CFNSD0 ) ,.FSWS8 ( FSWS8 )
     ,.FSWS7 ( FSWS7 ) ,.FSWS6 ( FSWS6 ) ,.FSWS5 ( FSWS5 ) ,.FSWS4 ( FSWS4 )
     ,.FSWS3 ( FSWS3 ) ,.FSWS2 ( FSWS2 ) ,.FSWS1 ( FSWS1 ) ,.FSWS0 ( FSWS0 )
     ,.FSWE9 ( FSWE9 ) ,.FSWE8 ( FSWE8 ) ,.FSWE7 ( FSWE7 ) ,.FSWE6 ( FSWE6 )
     ,.FSWE5 ( FSWE5 ) ,.FSWE4 ( FSWE4 ) ,.FSWE3 ( FSWE3 ) ,.FSWE2 ( FSWE2 )
     ,.FSWE1 ( FSWE1 ) ,.FSWE0 ( FSWE0 ) ,.CSPDTFLG ( CSPDTFLG ) ,.PBRAMEN ( pull_up49 )
     ,.SCANMODE ( SCANMODE ) ,.SCANRESZ ( SCANRESZ ) ,.PRDATA15 ( PRDMAW15 )
     ,.PRDATA14 ( PRDMAW14 ) ,.PRDATA13 ( PRDMAW13 ) ,.PRDATA12 ( PRDMAW12 )
     ,.PRDATA11 ( PRDMAW11 ) ,.PRDATA10 ( PRDMAW10 ) ,.PRDATA9 ( PRDMAW9 )
     ,.PRDATA8 ( PRDMAW8 ) ,.PRDATA7 ( PRDMAW7 ) ,.PRDATA6 ( PRDMAW6 )
     ,.PRDATA5 ( PRDMAW5 ) ,.PRDATA4 ( PRDMAW4 ) ,.PRDATA3 ( PRDMAW3 )
     ,.PRDATA2 ( PRDMAW2 ) ,.PRDATA1 ( PRDMAW1 ) ,.PRDATA0 ( PRDMAW0 )
     ,.DETECT ( DETECT ) ,.ICESVSTOP ( ICESVSTOP ) ,.ICEFETCHFLT ( ICEFETCHFLT )
     ,.ICEDATAFLT ( ICEDATAFLT ) ,.ICEDMAFLT ( ICEDMAFLT ) ,.ICECK60M ( ICECK60M )
    
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/_ice/_macro/_sss/modectl/100729/qlk0rmodectl2v1.hdl_nosec
  QLK0RMODECTL2V1 modectl (
    .POCRELNF ( POCRELNF ) ,.TRESET ( TRESET ) ,.RESETB ( RESETB ) ,.RESB ( RESB )
     ,.NSRESB ( NSRESB ) ,.PERESETZ ( RESB ) ,.RESETINBNF ( RESETINBNF )
     ,.BASECK ( BASECK ) ,.PCLKTST ( PCLKTST ) ,.TMDENCLK ( TMDENCLK )
     ,.BBMODE ( BBMODE ) ,.PRIMODIN ( HVIN ) ,.X2DIN ( X2DIN ) ,.C3HFF ( C3HFF )
     ,.SBRFONLY ( SBRFONLY ) ,.RXOCD ( RXOCD ) ,.UTI ( TIN00 ) ,.RNGIN6 ( pull_down15 )
     ,.RNGIN5 ( pull_down14 ) ,.RNGIN4 ( OSCOUTCP ) ,.RNGIN3 ( TFIHOCD )
     ,.RNGIN2 ( TFIHFL ) ,.RNGIN1 ( TR15KOUT ) ,.RNGIN0 ( TR32MOUT ) ,.ROUTSRC15 ( pull_down18 )
     ,.ROUTSRC14 ( pull_down17 ) ,.ROUTSRC13 ( DLY300NO ) ,.ROUTSRC12 ( P14EXINA )
     ,.ROUTSRC11 ( DLY50NO ) ,.ROUTSRC10 ( P13EXINA ) ,.ROUTSRC9 ( TLVIF )
     ,.ROUTSRC8 ( pull_down16 ) ,.ROUTSRC7 ( OSCOUTCP ) ,.ROUTSRC6 ( TFIHOCD )
     ,.ROUTSRC5 ( TFIHFL ) ,.ROUTSRC4 ( R15KSTPZ ) ,.ROUTSRC3 ( TR15KOUT )
     ,.ROUTSRC2 ( R32MSTP ) ,.ROUTSRC1 ( TR32MOUT ) ,.PSEL1 ( PSELMOD1 )
     ,.PSEL2 ( PSELMOD2 ) ,.PWRITE ( PWRITE ) ,.PENABLE ( PENABLE ) ,.GOFIRM ( GOFIRM )
     ,.PADDR1 ( PADDR1 ) ,.TESTMOD ( TESTMOD ) ,.FLMEMTES ( FLMEMTES )
     ,.SCANMODE ( SCANMODEICE ) ,.TESSCAN1 ( TESSCAN1 ) ,.TESSCAN2 ( TESSCAN2 )
     ,.TESSCAN3 ( TESSCAN3 ) ,.TESSCAN4 ( TESSCAN4 ) ,.TESINST ( TESINST )
     ,.BBTESINST ( BBTESINST ) ,.TESUSR ( TESUSR ) ,.TESDBT ( TESDBT )
     ,.TESTRMRD ( TESTRMRD ) ,.PTESINST ( PTESINST ) ,.OPTFLMEM ( OPTFLMEM )
     ,.OPTRAM ( OPTRAM ) ,.OPTIDDQ ( OPTIDDQ ) ,.PWDATA7 ( MDW7 ) ,.OPTEXCCK ( OPTEXCCK )
     ,.OPTOPLRD ( OPTOPLRD ) ,.OPTBCT ( OPTBCT ) ,.OPTDFL ( OPTDFL ) ,.OPTMDUMP ( OPTMDUMP )
     ,.RAMMULTI ( RAMMULTI ) ,.FMULTIEN ( FMULTIEN ) ,.MDLYCUT ( MDLYCUT )
     ,.RAEDIS ( RAEDIS ) ,.SLECCOFF ( SLECCOFF ) ,.SELTAR ( SELTAR ) ,.SELTAF ( SELTAF )
     ,.SELTADF ( SELTADF ) ,.PRDATA8 ( PRDMOD8 ) ,.STAYTES ( STAYTES )
     ,.TPIDSEL ( TPIDSEL ) ,.POSCOUTE ( POSCOUTE ) ,.POSCNOST ( POSCNOST )
     ,.OTI ( OTI00 ) ,.TESDBT2 ( TESDBT2 ) ,.GOFIRMR ( GOFIRMR ) ,.PADDR3 ( PADDR3 )
     ,.PADDR2 ( PADDR2 ) ,.PADDR0 ( PADDR0 ) ,.PWDATA15 ( MDW15 ) ,.PWDATA14 ( MDW14 )
     ,.PWDATA13 ( MDW13 ) ,.PWDATA12 ( MDW12 ) ,.PWDATA11 ( MDW11 ) ,.PWDATA10 ( MDW10 )
     ,.PWDATA9 ( MDW9 ) ,.PWDATA8 ( MDW8 ) ,.PWDATA6 ( MDW6 ) ,.PWDATA5 ( MDW5 )
     ,.PWDATA4 ( MDW4 ) ,.PWDATA3 ( MDW3 ) ,.PWDATA2 ( MDW2 ) ,.PWDATA1 ( MDW1 )
     ,.PWDATA0 ( MDW0 ) ,.PRDATA15 ( PRDMOD15 ) ,.PRDATA14 ( PRDMOD14 )
     ,.PRDATA13 ( PRDMOD13 ) ,.PRDATA12 ( PRDMOD12 ) ,.PRDATA11 ( PRDMOD11 )
     ,.PRDATA10 ( PRDMOD10 ) ,.PRDATA9 ( PRDMOD9 ) ,.PRDATA7 ( PRDMOD7 )
     ,.PRDATA6 ( PRDMOD6 ) ,.PRDATA5 ( PRDMOD5 ) ,.PRDATA4 ( PRDMOD4 )
     ,.PRDATA3 ( PRDMOD3 ) ,.PRDATA2 ( PRDMOD2 ) ,.PRDATA1 ( PRDMOD1 )
     ,.PRDATA0 ( PRDMOD0 ) ,.STBRELE ( STBRELE ) ,.HLTST ( HLTST ) ,.TID10 ( TID10 )
     ,.ECCER ( ECCER ) ,.DECCER ( DECCER ) ,.VCEQ ( VCEQ ) ,.RAMECCER ( pull_down13 )
     ,.MDR15 ( MDR15 ) ,.MDR14 ( MDR14 ) ,.MDR13 ( MDR13 ) ,.MDR12 ( MDR12 )
     ,.MDR11 ( MDR11 ) ,.MDR10 ( MDR10 ) ,.MDR9 ( MDR9 ) ,.MDR8 ( MDR8 )
     ,.MDR7 ( MDR7 ) ,.MDR6 ( MDR6 ) ,.MDR5 ( MDR5 ) ,.MDR4 ( MDR4 ) ,.MDR3 ( MDR3 )
     ,.MDR2 ( MDR2 ) ,.MDR1 ( MDR1 ) ,.MDR0 ( MDR0 ) ,.EIRAMO7 ( pull_down24 )
     ,.EIRAMO6 ( pull_down23 ) ,.EIRAMO5 ( pull_down22 ) ,.EIRAMO4 ( pull_down21 )
     ,.EIRAMO3 ( pull_down20 ) ,.EIRAMO2 ( pull_down19 ) ,.EIRAMO1 ( EIRAMO1 )
     ,.EIRAMO0 ( EIRAMO0 ) ,.RMULTIO23 ( pull_down48 ) ,.RMULTIO15 ( pull_down40 )
     ,.RMULTIO22 ( pull_down47 ) ,.RMULTIO14 ( pull_down39 ) ,.RMULTIO21 ( pull_down46 )
     ,.RMULTIO13 ( pull_down38 ) ,.RMULTIO20 ( pull_down45 ) ,.RMULTIO12 ( pull_down37 )
     ,.RMULTIO19 ( pull_down44 ) ,.RMULTIO18 ( pull_down43 ) ,.RMULTIO17 ( pull_down42 )
     ,.RMULTIO16 ( pull_down41 ) ,.RMULTIO11 ( pull_down36 ) ,.RMULTIO10 ( pull_down35 )
     ,.RMULTIO9 ( pull_down34 ) ,.RMULTIO8 ( pull_down33 ) ,.RMULTIO7 ( pull_down32 )
     ,.RMULTIO6 ( pull_down31 ) ,.RMULTIO5 ( pull_down30 ) ,.RMULTIO4 ( pull_down29 )
     ,.RMULTIO3 ( pull_down28 ) ,.RMULTIO2 ( pull_down27 ) ,.RMULTIO1 ( pull_down26 )
     ,.RMULTIO0 ( pull_down25 ) ,.FLRO37 ( FLRO37 ) ,.FLRO29 ( FLRO29 )
     ,.FLRO36 ( FLRO36 ) ,.FLRO28 ( FLRO28 ) ,.FLRO35 ( FLRO35 ) ,.FLRO27 ( FLRO27 )
     ,.FLRO19 ( FLRO19 ) ,.FLRO34 ( FLRO34 ) ,.FLRO26 ( FLRO26 ) ,.FLRO18 ( FLRO18 )
     ,.FLRO33 ( FLRO33 ) ,.FLRO25 ( FLRO25 ) ,.FLRO17 ( FLRO17 ) ,.FLRO32 ( FLRO32 )
     ,.FLRO24 ( FLRO24 ) ,.FLRO16 ( FLRO16 ) ,.FLRO31 ( FLRO31 ) ,.FLRO23 ( FLRO23 )
     ,.FLRO15 ( FLRO15 ) ,.FLRO30 ( FLRO30 ) ,.FLRO22 ( FLRO22 ) ,.FLRO14 ( FLRO14 )
     ,.FLRO21 ( FLRO21 ) ,.FLRO13 ( FLRO13 ) ,.FLRO20 ( FLRO20 ) ,.FLRO12 ( FLRO12 )
     ,.FLRO11 ( FLRO11 ) ,.FLRO10 ( FLRO10 ) ,.FLRO9 ( FLRO9 ) ,.FLRO8 ( FLRO8 )
     ,.FLRO7 ( FLRO7 ) ,.FLRO6 ( FLRO6 ) ,.FLRO5 ( FLRO5 ) ,.FLRO4 ( FLRO4 )
     ,.FLRO3 ( FLRO3 ) ,.FLRO2 ( FLRO2 ) ,.FLRO1 ( FLRO1 ) ,.FLRO0 ( FLRO0 )
     ,.DFLRO11 ( DFLRO11 ) ,.DFLRO10 ( DFLRO10 ) ,.DFLRO9 ( DFLRO9 ) ,.DFLRO8 ( DFLRO8 )
     ,.DFLRO7 ( DFLRO7 ) ,.DFLRO6 ( DFLRO6 ) ,.DFLRO5 ( DFLRO5 ) ,.DFLRO4 ( DFLRO4 )
     ,.DFLRO3 ( DFLRO3 ) ,.DFLRO2 ( DFLRO2 ) ,.DFLRO1 ( DFLRO1 ) ,.DFLRO0 ( DFLRO0 )
     ,.AF19 ( AF19 ) ,.AF18 ( AF18 ) ,.AF17 ( AF17 ) ,.AF16 ( AF16 ) ,.AF15 ( AF15 )
     ,.AF14 ( AF14 ) ,.AF13 ( AF13 ) ,.AF12 ( AF12 ) ,.AF11 ( AF11 ) ,.AF10 ( AF10 )
     ,.AF9 ( AF9 ) ,.AF8 ( AF8 ) ,.AF7 ( AF7 ) ,.AF6 ( AF6 ) ,.AF5 ( AF5 )
     ,.AF4 ( AF4 ) ,.AF3 ( AF3 ) ,.AF2 ( AF2 ) ,.CRCHLTEN ( CRCHLTEN )
     ,.INCDECMD ( INCDECMD ) ,.LFSSCAIN ( LFSSCAIN ) ,.MODERD ( MODERD )
     ,.MODEWR ( MODEWR ) ,.MODENOP ( MODENOP ) ,.MODEFNOP ( MODEFNOP )
     ,.INCDECWS1 ( INCDECWS1 ) ,.INCDECWS0 ( INCDECWS0 ) ,.TA17 ( TA17 )
     ,.TA16 ( TA16 ) ,.TA15 ( TA15 ) ,.TA14 ( TA14 ) ,.TA13 ( TA13 ) ,.TA12 ( TA12 )
     ,.TA11 ( TA11 ) ,.TA10 ( TA10 ) ,.TA9 ( TA9 ) ,.TA8 ( TA8 ) ,.TA7 ( TA7 )
     ,.TA6 ( TA6 ) ,.TA5 ( TA5 ) ,.TA4 ( TA4 ) ,.TA3 ( TA3 ) ,.TA2 ( TA2 )
     ,.TA1 ( TA1 ) ,.TA0 ( TA0 ) ,.SLFLASH ( SLFLASH ) ,.BTCLKIN ( R32MOUT )
     ,.RDSETUP ( RDSETUP ) ,.RESSQSTA ( RESSQSTA ) ,.RT0MON0 ( RT0MON0 )
     ,.RT0MON1 ( RT0MON1 ) ,.WDTMON ( WDTMON ) ,.SCANOUT ( pull_down52 )
     ,.TDIN5 ( TDIN5 ) ,.TDIN4 ( TDIN4 ) ,.TDIN3 ( TDIN3 ) ,.TDIN2T ( TDIN2T )
     ,.TDIN2R ( TDIN2R ) ,.TDIN1T ( TDIN1T ) ,.TDIN2B ( TDIN2B ) ,.TDIN2L ( pull_down49 )
     ,.TDIN1R ( TDIN1R ) ,.TDIN0T ( TDIN0T ) ,.TDIN1B ( TDIN1B ) ,.TDIN1L ( pull_down50 )
     ,.TDIN0R ( TDIN0R ) ,.TDIN0B ( TDIN0B ) ,.TDIN0L ( pull_down51 ) ,.WAITMOD ( WAITMOD )
     ,.EXCLK1 ( EXCLK1 ) ,.TID31 ( TID31 ) ,.TID23 ( TID23 ) ,.TID15 ( TID15 )
     ,.TID30 ( TID30 ) ,.TID22 ( TID22 ) ,.TID14 ( TID14 ) ,.TID29 ( TID29 )
     ,.TID28 ( TID28 ) ,.TID27 ( TID27 ) ,.TID19 ( TID19 ) ,.TID26 ( TID26 )
     ,.TID18 ( TID18 ) ,.TID25 ( TID25 ) ,.TID17 ( TID17 ) ,.TID24 ( TID24 )
     ,.TID16 ( TID16 ) ,.TID21 ( TID21 ) ,.TID13 ( TID13 ) ,.TID20 ( TID20 )
     ,.TID12 ( TID12 ) ,.TID11 ( TID11 ) ,.TID9 ( TID9 ) ,.TID8 ( TID8 )
     ,.TID7 ( TID7 ) ,.TID6 ( TID6 ) ,.TID5 ( TID5 ) ,.TID4 ( TID4 ) ,.TID3 ( TID3 )
     ,.TID2 ( TID2 ) ,.TID1 ( TID1 ) ,.TID0 ( TID0 ) ,.TESENI4 ( TESENI4 )
     ,.TESENI3 ( TESENI3 ) ,.TESENI2T ( TESENI2T ) ,.TESENI2R ( TESENI2R )
     ,.TESENI1T ( TESENI1T ) ,.TESENI2B ( TESENI2B ) ,.TESENI2L ( TESENI2L )
     ,.TESENI1R ( TESENI1R ) ,.TESENI0T ( TESENI0T ) ,.TESENI1B ( TESENI1B )
     ,.TESENI1L ( TESENI1L ) ,.TESENI0R ( TESENI0R ) ,.TESENI0B ( TESENI0B )
     ,.TESENI0L ( TESENI0L ) ,.TESENO3 ( TESENO3 ) ,.TESENO2T ( TESENO2T )
     ,.TESENO2R ( TESENO2R ) ,.TESENO1T ( TESENO1T ) ,.TESENO2B ( TESENO2B )
     ,.TESENO2L ( TESENO2L ) ,.TESENO1R ( TESENO1R ) ,.TESENO0T ( TESENO0T )
     ,.TESENO1B ( TESENO1B ) ,.TESENO1L ( TESENO1L ) ,.TESENO0R ( TESENO0R )
     ,.TESENO0B ( TESENO0B ) ,.TESENO0L ( TESENO0L ) ,.TDSEL3 ( TDSEL3 )
     ,.TDSEL2T ( TDSEL2T ) ,.TDSEL2R ( TDSEL2R ) ,.TDSEL1T ( TDSEL1T )
     ,.TDSEL2B ( TDSEL2B ) ,.TDSEL2L ( TDSEL2L ) ,.TDSEL1R ( TDSEL1R )
     ,.TDSEL0T ( TDSEL0T ) ,.TDSEL1B ( TDSEL1B ) ,.TDSEL1L ( TDSEL1L )
     ,.TDSEL0R ( TDSEL0R ) ,.TDSEL0B ( TDSEL0B ) ,.TDSEL0L ( TDSEL0L )
     ,.TDOUT3 ( TDOUT3 ) ,.TDOUT2 ( TDOUT2 ) ,.TDOUT1 ( TDOUT1 ) ,.TDOUT0 ( TDOUT0 )
     ,.SCANIN ( SCANIN ) ,.SCANCLK ( SCANCLKICE ) ,.SCANEN ( SCANENICE )
     ,.SCANRESZ ( SCANRESZICE ) ,.SCANENMD ( SCANENMD ) ,.TIIDER ( TIIDER )
     ,.BBSCANOUT ( BBSCANOUT )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/_ice/_macro/_sss/scon/100910/qlk0rscon1v1.hdl
  QLK0RSCON1V1 scon (
    .RESETB ( RESETB ) ,.SYSRESB ( SYSRESB ) ,.BASECK ( BASECK ) ,.TESINST ( TESINST )
     ,.CSPDTFLG ( CSPDTFLG ) ,.SVSTOP ( SVSTOP ) ,.PENABLE ( PENABLE )
     ,.PSEL ( PSELSCN ) ,.PADDR2 ( PADDR2 ) ,.PADDR1 ( PADDR1 ) ,.PADDR0 ( PADDR0 )
     ,.PWRITE ( PWRITE ) ,.SCANMODE ( SCANMODE ) ,.SCANRESZ ( SCANRESZ )
     ,.PRDATA15 ( PRDSCN15 ) ,.PRDATA14 ( PRDSCN14 ) ,.PRDATA13 ( PRDSCN13 )
     ,.PRDATA12 ( PRDSCN12 ) ,.PRDATA11 ( PRDSCN11 ) ,.PRDATA10 ( PRDSCN10 )
     ,.PRDATA9 ( PRDSCN9 ) ,.PRDATA8 ( PRDSCN8 ) ,.PRDATA7 ( PRDSCN7 )
     ,.PRDATA6 ( PRDSCN6 ) ,.PRDATA5 ( PRDSCN5 ) ,.PRDATA4 ( PRDSCN4 )
     ,.PRDATA3 ( PRDSCN3 ) ,.PRDATA2 ( PRDSCN2 ) ,.PRDATA1 ( PRDSCN1 )
     ,.PRDATA0 ( PRDSCN0 ) ,.SRESIN3 ( pull_down53 ) ,.SRESIN2 ( DETECT )
     ,.SRESIN1 ( ICECKSMER ) ,.SRESIN0 ( PSEUDOTIIDER ) ,.SFRESEN3 ( pull_down55 )
     ,.SFRESEN2 ( pull_up59 ) ,.SFRESEN1 ( pull_up58 ) ,.SFRESEN0 ( pull_down54 )
     ,.SRESREQ ( SRESREQ ) ,.PWDATA7 ( MDW7 ) ,.BBTESINST ( BBTESINST )
     ,.ICECK60M ( ICECK60M )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_2.0/_macro/_local/_timing_fix_macro/kx4_flashclk_dly_mf3_v1.00/kx4_flashclk_dly.hdl
  KX4_FLASHCLK_DLY flashclk_dly (
    .RDCLKC1 ( RDCLKC1 ) ,.BASECKHS ( BASECKHS )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/qnsc3ncp1v2_mf3_CF1.3_20100903-01/_misc/lib/MF3/cmos1_2.1V/verilog/QNSC3NCP1V2.v
  QNSC3NCP1V2 flash_cp (
    .BG1ST ( BG1ST ) ,.HVPPTS1 ( HVPPTS1 ) ,.FLREGENB ( FLREGENB ) ,.OSCOUT ( OSCOUTCP )
     ,.REQFL ( REQFL ) ,.RDSETUP ( RDSETUP ) ,.REG125ST ( REG125ST ) ,.SRCUT ( SRCUT )
     ,.SRCUTCP ( SRCUTCP ) ,.TRMRD1 ( TRMRD1 ) ,.TRMRD2 ( TRMRD2 ) ,.TRMRD1CK ( TRMRD1CK )
     ,.TRMRD2CK ( TRMRD2CK ) ,.VBRESZCP ( VBRESZCP ) ,.VCPHV ( VCPHV )
     ,.VPBIAS ( VPBIAS ) ,.VREGMV ( VREGMV ) ,.VREGRMV ( VREGRMV ) ,.VPPTS1 ( VPPTS1_CP )
     ,.CE ( CE0 ) ,.CER ( CER ) ,.CLKSEL1 ( CLKSEL1 ) ,.CPBT ( CPBT ) ,.CPT ( CPT )
     ,.CWEE ( CWEE ) ,.DCE ( DCE0 ) ,.DCER ( DCER ) ,.DCLKSEL1 ( DCLKSEL1 )
     ,.DDIS ( DDIS ) ,.DFLSTOP ( DFLSTOP ) ,.DIS ( DIS ) ,.DMRG00 ( DMRG00 )
     ,.DMRG01 ( DMRG01 ) ,.DMRG10 ( DMRG10 ) ,.DMRG11 ( DMRG11 ) ,.DMRG12 ( DMRG12 )
     ,.DRDCLKC1 ( DRDCLKC1 ) ,.DREAD ( DREAD ) ,.DSER ( DSER ) ,.DWED ( DWED )
     ,.DWWR ( DWWR ) ,.EXER ( EXER ) ,.EXTVPP1 ( EXTVPP1 ) ,.EXTVPP2 ( EXTVPP2 )
     ,.FCLK1 ( FCLK1 ) ,.FLSTOP ( FLSTOP ) ,.HISPEED ( HISPEED ) ,.IONCHK1 ( IONCHK1 )
     ,.IREFT ( IREFT ) ,.LOWPOWER ( LOWPOWER ) ,.LOWSPY ( LOWSPY ) ,.MEOC ( MEOC )
     ,.MEOR ( MEOR ) ,.MRG00 ( MRG00 ) ,.MRG01 ( MRG01 ) ,.MRG10 ( MRG10 )
     ,.MRG11 ( MRG11 ) ,.MRG12 ( MRG12 ) ,.MSWR ( MSWR ) ,.OSCNOSTP ( OSCNOSTP )
     ,.OSCOUTEN ( OSCOUTEN ) ,.POCREL ( POCRELNF ) ,.PROGI ( PROGI ) ,.RDCLKC1 ( RDCLKC1 )
     ,.RDCLKP1 ( RDCLKP1 ) ,.RDMRG0 ( RDMRG0 ) ,.RDMRG1 ( RDMRG1 ) ,.RDMRGC ( RDMRGC )
     ,.FIHFL ( FIHFL ) ,.RDT ( RDT ) ,.READ ( READ ) ,.POCREL5V ( POCREL5V )
     ,.RLOWSPY ( RLOWSPY ) ,.RTRMCP15 ( RTRMCP015 ) ,.RTRMCP16 ( RTRMCP016 )
     ,.RTRMCP17 ( RTRMCP017 ) ,.RTRMCP18 ( RTRMCP018 ) ,.RTRMCP19 ( RTRMCP019 )
     ,.RTRMCP20 ( RTRMCP020 ) ,.SCANMODE ( SCANMODE ) ,.SER ( SER ) ,.STCHK ( STCHK )
     ,.SUB ( SUB ) ,.TESDBT ( TESDBT ) ,.TRMCP0 ( TRMCP00 ) ,.TRMCP1 ( TRMCP01 )
     ,.TRMCP2 ( TRMCP02 ) ,.TRMCP3 ( TRMCP03 ) ,.TRMCP4 ( TRMCP04 ) ,.TRMCP5 ( TRMCP05 )
     ,.TRMCP6 ( TRMCP06 ) ,.TRMCP7 ( TRMCP07 ) ,.TRMCP8 ( TRMCP08 ) ,.TRMCP9 ( TRMCP09 )
     ,.TRMCP15 ( TRMCP015 ) ,.TRMCP16 ( TRMCP016 ) ,.TRMCP17 ( TRMCP017 )
     ,.VBRESZ ( RESETB ) ,.VREG ( VREG ) ,.WDT1 ( WDT1 ) ,.WDT2 ( WDT2 )
     ,.WDT3 ( WDT3 ) ,.WDT4 ( WDT4 ) ,.WED ( WED ) ,.WWR ( WWR ) ,.VCPRGWE ( VCPRGWE )
     ,.RESB ( RESB )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/qnsc3nreg1v2_mf3_CF1.3_20100903-01/_misc/lib/MF3/cmos1_2.1V/verilog/QNSC3NREG1V2.v
  QNSC3NREG1V2 flash_reg (
    .POCREL5V ( POCREL5V ) ,.FLREGENB ( FLREGENB ) ,.VCPRGWE ( VCPRGWE )
    
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/qnsc3ncpdc0v1_mf3_CF1.3_20100903-01/_misc/lib/MF3/cmos1_2.1V/verilog/QNSC3NCPDC0V1.v
  QNSC3NCPDC0V1 flash_capa0 (
    .VCPHV ( VCPHV )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/qnsc3ncpdc0v1_mf3_CF1.3_20100903-01/_misc/lib/MF3/cmos1_2.1V/verilog/QNSC3NCPDC0V1.v
  QNSC3NCPDC0V1 flash_capa1 (
    .VCPHV ( VCPHV )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/qnsc3ncpdc0v1_mf3_CF1.3_20100903-01/_misc/lib/MF3/cmos1_2.1V/verilog/QNSC3NCPDC0V1.v
  QNSC3NCPDC0V1 flash_capa2 (
    .VCPHV ( VCPHV )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/qnsc3ncpdc0v1_mf3_CF1.3_20100903-01/_misc/lib/MF3/cmos1_2.1V/verilog/QNSC3NCPDC0V1.v
  QNSC3NCPDC0V1 flash_capa3 (
    .VCPHV ( VCPHV )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/qnsc3ncpdc0v1_mf3_CF1.3_20100903-01/_misc/lib/MF3/cmos1_2.1V/verilog/QNSC3NCPDC0V1.v
  QNSC3NCPDC0V1 flash_capa4 (
    .VCPHV ( VCPHV )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/qnsc3ncpdc0v1_mf3_CF1.3_20100903-01/_misc/lib/MF3/cmos1_2.1V/verilog/QNSC3NCPDC0V1.v
  QNSC3NCPDC0V1 flash_capa5 (
    .VCPHV ( VCPHV )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/qnsc3ncpdc0v1_mf3_CF1.3_20100903-01/_misc/lib/MF3/cmos1_2.1V/verilog/QNSC3NCPDC0V1.v
  QNSC3NCPDC0V1 flash_capa6 (
    .VCPHV ( VCPHV )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/qnsc3ncpdc0v1_mf3_CF1.3_20100903-01/_misc/lib/MF3/cmos1_2.1V/verilog/QNSC3NCPDC0V1.v
  QNSC3NCPDC0V1 flash_capa7 (
    .VCPHV ( VCPHV )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/qnsc3ncpdc0v1_mf3_CF1.3_20100903-01/_misc/lib/MF3/cmos1_2.1V/verilog/QNSC3NCPDC0V1.v
  QNSC3NCPDC0V1 flash_capa8 (
    .VCPHV ( VCPHV )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/qnsc3ncpdc0v1_mf3_CF1.3_20100903-01/_misc/lib/MF3/cmos1_2.1V/verilog/QNSC3NCPDC0V1.v
  QNSC3NCPDC0V1 flash_capa9 (
    .VCPHV ( VCPHV )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/qnsc3ncpdc0v1_mf3_CF1.3_20100903-01/_misc/lib/MF3/cmos1_2.1V/verilog/QNSC3NCPDC0V1.v
  QNSC3NCPDC0V1 flash_capa10 (
    .VCPHV ( VCPHV )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/qnsc3ncpdc0v1_mf3_CF1.3_20100903-01/_misc/lib/MF3/cmos1_2.1V/verilog/QNSC3NCPDC0V1.v
  QNSC3NCPDC0V1 flash_capa11 (
    .VCPHV ( VCPHV )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/qnsc3ncpdc0v1_mf3_CF1.3_20100903-01/_misc/lib/MF3/cmos1_2.1V/verilog/QNSC3NCPDC0V1.v
  QNSC3NCPDC0V1 flash_capa12 (
    .VCPHV ( VCPHV )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/qnsc3ncpdc0v1_mf3_CF1.3_20100903-01/_misc/lib/MF3/cmos1_2.1V/verilog/QNSC3NCPDC0V1.v
  QNSC3NCPDC0V1 flash_capa13 (
    .VCPHV ( VCPHV )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/qnsc3ncpdc0v1_mf3_CF1.3_20100903-01/_misc/lib/MF3/cmos1_2.1V/verilog/QNSC3NCPDC0V1.v
  QNSC3NCPDC0V1 flash_capa14 (
    .VCPHV ( VCPHV )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_2.0/_macro/_local/kx4_busbridge_mf3_v2.00/_library/100821/kx4_busbridge.hdl
  KX4_BUSBRIDGE bbr (
    .SLMEM ( SLMEM ) ,.CPURD ( CPURD ) ,.CPUWR ( CPUWR ) ,.MA15 ( MA15 )
     ,.MA14 ( MA14 ) ,.MA13 ( MA13 ) ,.MA12 ( MA12 ) ,.MA11 ( MA11 ) ,.MA10 ( MA10 )
     ,.MA9 ( MA9 ) ,.MA8 ( MA8 ) ,.MA7 ( MA7 ) ,.MA6 ( MA6 ) ,.MA5 ( MA5 )
     ,.MA4 ( MA4 ) ,.MA3 ( MA3 ) ,.MA2 ( MA2 ) ,.MA1 ( MA1 ) ,.MA0 ( MA0 )
     ,.MDW15 ( MDW15 ) ,.MDW14 ( MDW14 ) ,.MDW13 ( MDW13 ) ,.MDW12 ( MDW12 )
     ,.MDW11 ( MDW11 ) ,.FLRO9 ( FLRO9 ) ,.MDW10 ( MDW10 ) ,.FLRO8 ( FLRO8 )
     ,.MDW9 ( MDW9 ) ,.MDW8 ( MDW8 ) ,.MDW7 ( MDW7 ) ,.MDW6 ( MDW6 ) ,.MDW5 ( MDW5 )
     ,.MDW4 ( MDW4 ) ,.MDW3 ( MDW3 ) ,.MDW2 ( MDW2 ) ,.MDW1 ( MDW1 ) ,.MDW0 ( MDW0 )
     ,.BBMODE ( BBMODE ) ,.BBNVM1 ( BBNVM1 ) ,.BBNVM2 ( BBNVM2 ) ,.BBTESINST ( BBTESINST )
     ,.PRDSELEN ( PRDSELEN ) ,.PRDRTC12 ( PRDRTC12 ) ,.FLRO15 ( FLRO15 )
     ,.FLRO14 ( FLRO14 ) ,.FLRO13 ( FLRO13 ) ,.FLRO12 ( FLRO12 ) ,.FLRO11 ( FLRO11 )
     ,.FLRO10 ( FLRO10 ) ,.FLRO7 ( FLRO7 ) ,.FLRO6 ( FLRO6 ) ,.FLRO5 ( FLRO5 )
     ,.FLRO4 ( FLRO4 ) ,.FLRO3 ( FLRO3 ) ,.FLRO2 ( FLRO2 ) ,.FLRO1 ( FLRO1 )
     ,.FLRO0 ( FLRO0 ) ,.MDRRAM15 ( MDRRAM15 ) ,.MDRRAM14 ( MDRRAM14 )
     ,.MDRRAM13 ( MDRRAM13 ) ,.MDRRAM12 ( MDRRAM12 ) ,.MDRRAM11 ( MDRRAM11 )
     ,.MDRRAM10 ( MDRRAM10 ) ,.MDRRAM9 ( MDRRAM9 ) ,.MDRRAM8 ( MDRRAM8 )
     ,.MDRRAM7 ( MDRRAM7 ) ,.MDRRAM6 ( MDRRAM6 ) ,.MDRRAM5 ( MDRRAM5 )
     ,.MDRRAM4 ( MDRRAM4 ) ,.MDRRAM3 ( MDRRAM3 ) ,.MDRINT9 ( MDRINT9 )
     ,.MDRRAM2 ( MDRRAM2 ) ,.MDRINT8 ( MDRINT8 ) ,.MDRRAM1 ( MDRRAM1 )
     ,.MDRINT7 ( MDRINT7 ) ,.MDRRAM0 ( MDRRAM0 ) ,.MDRINT6 ( MDRINT6 )
     ,.MDRMUL15 ( MDRMUL15 ) ,.MDRMUL14 ( MDRMUL14 ) ,.MDRMUL13 ( MDRMUL13 )
     ,.MDRMUL12 ( MDRMUL12 ) ,.MDRMUL11 ( MDRMUL11 ) ,.MDRMUL10 ( MDRMUL10 )
     ,.MDRMUL9 ( MDRMUL9 ) ,.PENABLE ( PENABLE ) ,.MDRMUL8 ( MDRMUL8 )
     ,.MDRMUL7 ( MDRMUL7 ) ,.MDRMUL6 ( MDRMUL6 ) ,.MDRMUL5 ( MDRMUL5 )
     ,.MDRMUL4 ( MDRMUL4 ) ,.MDRMUL3 ( MDRMUL3 ) ,.MDRMUL2 ( MDRMUL2 )
     ,.MDRMUL1 ( MDRMUL1 ) ,.MDRMUL0 ( MDRMUL0 ) ,.MDRINT15 ( MDRINT15 )
     ,.MDRINT14 ( MDRINT14 ) ,.MDRINT13 ( MDRINT13 ) ,.MDRINT12 ( MDRINT12 )
     ,.MDRINT11 ( MDRINT11 ) ,.MDRINT10 ( MDRINT10 ) ,.MDRINT5 ( MDRINT5 )
     ,.MDRINT4 ( MDRINT4 ) ,.MDRINT3 ( MDRINT3 ) ,.MDRINT2 ( MDRINT2 )
     ,.MDRINT1 ( MDRINT1 ) ,.MDRINT0 ( MDRINT0 ) ,.MDRDMA15 ( MDRDMA15 )
     ,.MDRDMA14 ( MDRDMA14 ) ,.MDRDMA13 ( MDRDMA13 ) ,.MDRDMA12 ( MDRDMA12 )
     ,.MDRDMA11 ( MDRDMA11 ) ,.MDRDMA10 ( MDRDMA10 ) ,.MDRDMA9 ( MDRDMA9 )
     ,.MDRDMA8 ( MDRDMA8 ) ,.MDRDMA7 ( MDRDMA7 ) ,.MDRDMA6 ( MDRDMA6 )
     ,.MDRDMA5 ( MDRDMA5 ) ,.MDRDMA4 ( MDRDMA4 ) ,.MDRDMA3 ( MDRDMA3 )
     ,.MDRDMA2 ( MDRDMA2 ) ,.MDRDMA1 ( MDRDMA1 ) ,.MDRDMA0 ( MDRDMA0 )
     ,.MDROCD15 ( MDROCD15 ) ,.MDROCD14 ( MDROCD14 ) ,.MDROCD13 ( MDROCD13 )
     ,.MDROCD12 ( MDROCD12 ) ,.MDROCD11 ( MDROCD11 ) ,.MDROCD10 ( MDROCD10 )
     ,.MDROCD9 ( MDROCD9 ) ,.MDROCD8 ( MDROCD8 ) ,.MDROCD7 ( MDROCD7 )
     ,.MDROCD6 ( MDROCD6 ) ,.MDROCD5 ( MDROCD5 ) ,.MDROCD4 ( MDROCD4 )
     ,.MDROCD3 ( MDROCD3 ) ,.MDROCD2 ( MDROCD2 ) ,.MDROCD1 ( MDROCD1 )
     ,.MDROCD0 ( MDROCD0 ) ,.MDRIM815 ( MDRIM815 ) ,.MDRIM814 ( MDRIM814 )
     ,.MDRIM813 ( MDRIM813 ) ,.MDRIM812 ( MDRIM812 ) ,.MDRIM811 ( MDRIM811 )
     ,.MDRIM810 ( MDRIM810 ) ,.MDRIM89 ( MDRIM89 ) ,.MDRIM88 ( MDRIM88 )
     ,.MDRIM87 ( MDRIM87 ) ,.MDRIM86 ( MDRIM86 ) ,.MDRIM85 ( MDRIM85 )
     ,.MDRIM84 ( MDRIM84 ) ,.MDRIM83 ( MDRIM83 ) ,.MDRIM82 ( MDRIM82 )
     ,.MDRIM81 ( MDRIM81 ) ,.MDRIM49 ( MDRIM49 ) ,.MDRIM80 ( MDRIM80 )
     ,.MDRIM48 ( MDRIM48 ) ,.MDRIM411 ( MDRIM411 ) ,.MDRIM410 ( MDRIM410 )
     ,.MDRIM43 ( MDRIM43 ) ,.MDRIM42 ( MDRIM42 ) ,.MDRIM41 ( MDRIM41 )
     ,.MDRIM40 ( MDRIM40 ) ,.MDRPOG15 ( MDRPOG15 ) ,.MDRPOG14 ( MDRPOG14 )
     ,.MDRPOG13 ( MDRPOG13 ) ,.MDRPOG12 ( MDRPOG12 ) ,.MDRPOG11 ( MDRPOG11 )
     ,.MDRPOG10 ( MDRPOG10 ) ,.MDRPOG9 ( MDRPOG9 ) ,.MDRPOG8 ( MDRPOG8 )
     ,.MDRPOG7 ( MDRPOG7 ) ,.MDRPOG6 ( MDRPOG6 ) ,.MDRPOG5 ( MDRPOG5 )
     ,.MDRPOG4 ( MDRPOG4 ) ,.MDRPOG3 ( MDRPOG3 ) ,.MDRPOG2 ( MDRPOG2 )
     ,.MDRPOG1 ( MDRPOG1 ) ,.MDRPOG0 ( MDRPOG0 ) ,.MDRCID15 ( MDRCID15 )
     ,.MDRCID14 ( MDRCID14 ) ,.MDRCID13 ( MDRCID13 ) ,.MDRCID12 ( MDRCID12 )
     ,.MDRCID11 ( MDRCID11 ) ,.MDRCID10 ( MDRCID10 ) ,.MDRCID9 ( MDRCID9 )
     ,.MDRCID8 ( MDRCID8 ) ,.MDRCID7 ( MDRCID7 ) ,.MDRCID6 ( MDRCID6 )
     ,.MDRCID5 ( MDRCID5 ) ,.MDRCID4 ( MDRCID4 ) ,.MDRCID3 ( MDRCID3 )
     ,.MDRCID2 ( MDRCID2 ) ,.MDRCID1 ( MDRCID1 ) ,.MDRCID0 ( MDRCID0 )
     ,.PRDCSC15 ( PRDCSC15 ) ,.PRDCSC14 ( PRDCSC14 ) ,.PRDCSC13 ( PRDCSC13 )
     ,.PRDCSC12 ( PRDCSC12 ) ,.PRDCSC11 ( PRDCSC11 ) ,.PRDCSC10 ( PRDCSC10 )
     ,.PRDCSC9 ( PRDCSC9 ) ,.PRDIIC1 ( PRDIIC1 ) ,.PRDCSC8 ( PRDCSC8 )
     ,.PRDIIC0 ( PRDIIC0 ) ,.PRDCSC7 ( PRDCSC7 ) ,.PRDCSC6 ( PRDCSC6 )
     ,.PRDCSC5 ( PRDCSC5 ) ,.PRDCRC9 ( PRDCRC9 ) ,.PRDCSC4 ( PRDCSC4 )
     ,.PRDCRC8 ( PRDCRC8 ) ,.PRDCSC3 ( PRDCSC3 ) ,.PRDCRC7 ( PRDCRC7 )
     ,.PRDCSC2 ( PRDCSC2 ) ,.PRDCRC6 ( PRDCRC6 ) ,.PRDCSC1 ( PRDCSC1 )
     ,.PRDCRC5 ( PRDCRC5 ) ,.PRDCSC0 ( PRDCSC0 ) ,.PRDCRC4 ( PRDCRC4 )
     ,.PRDPCL15 ( PRDPCL15 ) ,.PRDPCL14 ( pull_down56 ) ,.PRDPCL13 ( pull_down57 )
     ,.PRDPCL12 ( pull_down58 ) ,.PRDPCL11 ( PRDPCL11 ) ,.PRDPCL10 ( PRDPCL10 )
     ,.PRDPCL9 ( PRDPCL9 ) ,.PRDMOD1 ( PRDMOD1 ) ,.PRDPCL8 ( PRDPCL8 )
     ,.PRDMOD0 ( PRDMOD0 ) ,.PRDPCL7 ( PRDPCL7 ) ,.PRDPCL6 ( pull_down59 )
     ,.PRDPCL5 ( pull_down60 ) ,.PRDPCL4 ( pull_down61 ) ,.PRDPCL3 ( PRDPCL3 )
     ,.PRDPCL2 ( PRDPCL2 ) ,.PRDPCL1 ( PRDPCL1 ) ,.PRDPCL0 ( PRDPCL0 )
     ,.PRDMOD15 ( PRDMOD15 ) ,.PRDMOD14 ( PRDMOD14 ) ,.PRDMOD13 ( PRDMOD13 )
     ,.PRDMOD12 ( PRDMOD12 ) ,.PRDMOD11 ( PRDMOD11 ) ,.PRDMOD10 ( PRDMOD10 )
     ,.PRDMOD9 ( PRDMOD9 ) ,.PSELP13 ( PSELP13 ) ,.PRDMOD8 ( PRDMOD8 )
     ,.PSELP12 ( PSELP12 ) ,.PRDMOD7 ( PRDMOD7 ) ,.PRDMOD6 ( PRDMOD6 )
     ,.PSELBCD ( PSELBCD ) ,.PRDMOD5 ( PRDMOD5 ) ,.PRDMOD4 ( PRDMOD4 )
     ,.PRDMOD3 ( PRDMOD3 ) ,.PRDMOD2 ( PRDMOD2 ) ,.PRDWDT15 ( PRDWDT15 )
     ,.PRDWDT12 ( PRDWDT12 ) ,.PRDWDT11 ( PRDWDT11 ) ,.PRDWDT9 ( PRDWDT9 )
     ,.PRDFCB15 ( PRDFCB15 ) ,.PRDCIC11 ( PRDCIC11 ) ,.PRDFCB14 ( PRDFCB14 )
     ,.PRDCIC10 ( PRDCIC10 ) ,.PRDFCB13 ( PRDFCB13 ) ,.PRDFCB12 ( PRDFCB12 )
     ,.PRDFCB11 ( PRDFCB11 ) ,.PRDFCB10 ( PRDFCB10 ) ,.PRDFCB9 ( PRDFCB9 )
     ,.PRDCIC7 ( PRDCIC7 ) ,.PRDCID5 ( PRDCID5 ) ,.PRDFCB8 ( PRDFCB8 )
     ,.PRDCIC6 ( PRDCIC6 ) ,.PRDCID4 ( PRDCID4 ) ,.PRDFCB7 ( PRDFCB7 )
     ,.PRDCIC5 ( PRDCIC5 ) ,.PRDCID3 ( PRDCID3 ) ,.PRDFCB6 ( PRDFCB6 )
     ,.PRDCIC4 ( PRDCIC4 ) ,.PRDCID2 ( PRDCID2 ) ,.PRDFCB5 ( PRDFCB5 )
     ,.PRDCIC3 ( PRDCIC3 ) ,.PRDCID1 ( PRDCID1 ) ,.PRDFCB4 ( PRDFCB4 )
     ,.PRDCIC2 ( PRDCIC2 ) ,.PRDCID0 ( PRDCID0 ) ,.PRDFCB3 ( PRDFCB3 )
     ,.PRDCIC1 ( PRDCIC1 ) ,.PRDFCB2 ( PRDFCB2 ) ,.PRDCIC0 ( PRDCIC0 )
     ,.PRDFCB1 ( PRDFCB1 ) ,.PRDFCB0 ( PRDFCB0 ) ,.PRDRTC15 ( PRDRTC15 )
     ,.PRDRTC14 ( PRDRTC14 ) ,.PRDRTC13 ( PRDRTC13 ) ,.PRDRTC11 ( PRDRTC11 )
     ,.PRDRTC10 ( PRDRTC10 ) ,.PSELOCD2 ( PSELOCD2 ) ,.PRDRTC9 ( PRDRTC9 )
     ,.PRDRTC8 ( PRDRTC8 ) ,.PRDRTC7 ( PRDRTC7 ) ,.PSELMAW ( PSELMAW )
     ,.PRDRTC6 ( PRDRTC6 ) ,.PRDRTC5 ( PRDRTC5 ) ,.WAITMEM ( WAITMEM )
     ,.PRDRTC4 ( PRDRTC4 ) ,.PRDRTC3 ( PRDRTC3 ) ,.PRDRTC2 ( PRDRTC2 )
     ,.PRDRTC1 ( PRDRTC1 ) ,.PRDRTC0 ( PRDRTC0 ) ,.PRDIIC15 ( PRDIIC15 )
     ,.PRDIIC14 ( PRDIIC14 ) ,.PRDIIC13 ( PRDIIC13 ) ,.PRDIIC12 ( PRDIIC12 )
     ,.PRDIIC11 ( PRDIIC11 ) ,.PRDIIC10 ( PRDIIC10 ) ,.PRDIIC9 ( PRDIIC9 )
     ,.PRDIIC8 ( PRDIIC8 ) ,.PRDIIC7 ( PRDIIC7 ) ,.PRDIIC6 ( PRDIIC6 )
     ,.PRDIIC5 ( PRDIIC5 ) ,.PRDIIC4 ( PRDIIC4 ) ,.PRDIIC3 ( PRDIIC3 )
     ,.PRDIIC2 ( PRDIIC2 ) ,.PRDTA015 ( PRDTA015 ) ,.PRDTA014 ( PRDTA014 )
     ,.PRDTA013 ( PRDTA013 ) ,.PRDTA012 ( PRDTA012 ) ,.PRDTA011 ( PRDTA011 )
     ,.PRDTA010 ( PRDTA010 ) ,.PRDTA09 ( PRDTA09 ) ,.PRDTA08 ( PRDTA08 )
     ,.PRDTA07 ( PRDTA07 ) ,.PRDTA06 ( PRDTA06 ) ,.PRDTA05 ( PRDTA05 )
     ,.PRDTA04 ( PRDTA04 ) ,.PRDTA03 ( PRDTA03 ) ,.PRDSA19 ( PRDSA19 )
     ,.PRDTA02 ( PRDTA02 ) ,.PRDSA18 ( PRDSA18 ) ,.PRDTA01 ( PRDTA01 )
     ,.PRDSA09 ( PRDSA09 ) ,.PRDSA17 ( PRDSA17 ) ,.PRDTA00 ( PRDTA00 )
     ,.PRDSA08 ( PRDSA08 ) ,.PRDSA16 ( PRDSA16 ) ,.PRDSA015 ( PRDSA015 )
     ,.PRDSA111 ( PRDSA111 ) ,.PRDSA014 ( PRDSA014 ) ,.PRDSA110 ( PRDSA110 )
     ,.PRDSA013 ( PRDSA013 ) ,.PRDSA012 ( PRDSA012 ) ,.PRDSA011 ( PRDSA011 )
     ,.PRDSA010 ( PRDSA010 ) ,.PRDSA07 ( PRDSA07 ) ,.PRDSA15 ( PRDSA15 )
     ,.PRDSA06 ( PRDSA06 ) ,.PRDSA14 ( PRDSA14 ) ,.PRDSA05 ( PRDSA05 )
     ,.PRDSA13 ( PRDSA13 ) ,.PRDSA04 ( PRDSA04 ) ,.PRDSA12 ( PRDSA12 )
     ,.PRDSA03 ( PRDSA03 ) ,.PRDSA11 ( PRDSA11 ) ,.PRDSA02 ( PRDSA02 )
     ,.PRDSA10 ( PRDSA10 ) ,.PRDSA01 ( PRDSA01 ) ,.PRDSA00 ( PRDSA00 )
     ,.PRDSA115 ( PRDSA115 ) ,.PRDSA114 ( PRDSA114 ) ,.PRDSA113 ( PRDSA113 )
     ,.PRDSA112 ( PRDSA112 ) ,.PRDAD15 ( PRDAD15 ) ,.PRDAD14 ( PRDAD14 )
     ,.PRDAD13 ( PRDAD13 ) ,.PRDAD12 ( PRDAD12 ) ,.PRDAD11 ( PRDAD11 )
     ,.PRDAD10 ( PRDAD10 ) ,.PRDAD9 ( PRDAD9 ) ,.PRDAD8 ( PRDAD8 ) ,.PRDAD7 ( PRDAD7 )
     ,.PRDAD6 ( PRDAD6 ) ,.PRDAD5 ( PRDAD5 ) ,.PRDAD4 ( PRDAD4 ) ,.PRDAD3 ( PRDAD3 )
     ,.PRDAD2 ( PRDAD2 ) ,.PRDAD1 ( PRDAD1 ) ,.PRDAD0 ( PRDAD0 ) ,.PRDCIC15 ( PRDCIC15 )
     ,.PRDCID11 ( PRDCID11 ) ,.PRDCIC14 ( PRDCIC14 ) ,.PRDCID10 ( PRDCID10 )
     ,.PRDCIC13 ( PRDCIC13 ) ,.PRDCIC12 ( PRDCIC12 ) ,.PRDCIC9 ( PRDCIC9 )
     ,.PRDCID7 ( PRDCID7 ) ,.PRDCIC8 ( PRDCIC8 ) ,.PRDCID6 ( PRDCID6 )
     ,.PRDCID15 ( PRDCID15 ) ,.PRDCID14 ( PRDCID14 ) ,.PRDCID13 ( PRDCID13 )
     ,.PRDCID12 ( PRDCID12 ) ,.PRDCID9 ( PRDCID9 ) ,.PRDCID8 ( PRDCID8 )
     ,.PRDP0007 ( PRDP0007 ) ,.PRDP0111 ( PRDP0111 ) ,.PRDP0006 ( PRDP0006 )
     ,.PRDP0110 ( PRDP0110 ) ,.PRDP0005 ( PRDP0005 ) ,.PRDP0004 ( PRDP0004 )
     ,.PRDP0003 ( PRDP0003 ) ,.PRDP0002 ( PRDP0002 ) ,.PRDP0001 ( PRDP0001 )
     ,.PRDP0000 ( PRDP0000 ) ,.PRDP0115 ( PRDP0115 ) ,.PRDP0203 ( PRDP0203 )
     ,.PRDP0114 ( PRDP0114 ) ,.PRDP0202 ( PRDP0202 ) ,.PRDP0113 ( PRDP0113 )
     ,.PRDP0201 ( PRDP0201 ) ,.PRDP0112 ( PRDP0112 ) ,.PRDP0200 ( PRDP0200 )
     ,.PRDP0109 ( PRDP0109 ) ,.PRDP0205 ( PRDP0205 ) ,.PRDP0108 ( PRDP0108 )
     ,.PRDP0204 ( PRDP0204 ) ,.PRDP0207 ( PRDP0207 ) ,.PRDP0311 ( PRDP0311 )
     ,.PRDP0206 ( PRDP0206 ) ,.PRDP0310 ( PRDP0310 ) ,.PRDP0315 ( PRDP0315 )
     ,.PRDP0403 ( PRDP0403 ) ,.PRDP1203 ( PRDP1203 ) ,.PRDP0314 ( PRDP0314 )
     ,.PRDP0402 ( PRDP0402 ) ,.PRDP1202 ( PRDP1202 ) ,.PRDP0313 ( PRDP0313 )
     ,.PRDP0401 ( PRDP0401 ) ,.PRDP1201 ( PRDP1201 ) ,.PRDP0312 ( PRDP0312 )
     ,.PRDP0400 ( PRDP0400 ) ,.PRDP1200 ( PRDP1200 ) ,.PRDP0309 ( PRDP0309 )
     ,.PRDP0405 ( PRDP0405 ) ,.PRDP1205 ( PRDP1205 ) ,.PRDP0308 ( PRDP0308 )
     ,.PRDP0404 ( PRDP0404 ) ,.PRDP1204 ( PRDP1204 ) ,.PRDP0407 ( PRDP0407 )
     ,.PRDP0511 ( PRDP0511 ) ,.PRDP1207 ( PRDP1207 ) ,.PRDP1311 ( PRDP1311 )
     ,.PRDP0406 ( PRDP0406 ) ,.PRDP0510 ( PRDP0510 ) ,.PRDP1206 ( PRDP1206 )
     ,.PRDP1310 ( PRDP1310 ) ,.PRDP0515 ( PRDP0515 ) ,.PRDP0603 ( PRDP0603 )
     ,.PRDP1315 ( PRDP1315 ) ,.PRDP1403 ( PRDP1403 ) ,.PRDP0514 ( PRDP0514 )
     ,.PRDP0602 ( PRDP0602 ) ,.PRDP1314 ( PRDP1314 ) ,.PRDP1402 ( PRDP1402 )
     ,.PRDP0513 ( PRDP0513 ) ,.PRDP0601 ( PRDP0601 ) ,.PRDP1313 ( PRDP1313 )
     ,.PRDP1401 ( PRDP1401 ) ,.PRDP0512 ( PRDP0512 ) ,.PRDP0600 ( PRDP0600 )
     ,.PRDP1312 ( PRDP1312 ) ,.PRDP1400 ( PRDP1400 ) ,.PRDP0509 ( PRDP0509 )
     ,.PRDP0605 ( PRDP0605 ) ,.PRDP1309 ( PRDP1309 ) ,.PRDP1405 ( PRDP1405 )
     ,.PRDP0508 ( PRDP0508 ) ,.PRDP0604 ( PRDP0604 ) ,.PRDP1308 ( PRDP1308 )
     ,.PRDP1404 ( PRDP1404 ) ,.PRDP0607 ( PRDP0607 ) ,.PRDP0711 ( PRDP0711 )
     ,.PRDP1407 ( PRDP1407 ) ,.PRDP0606 ( PRDP0606 ) ,.PRDP0710 ( PRDP0710 )
     ,.PRDP1406 ( PRDP1406 ) ,.PRDP0715 ( PRDP0715 ) ,.PRDP0714 ( PRDP0714 )
     ,.PRDP0713 ( PRDP0713 ) ,.PRDP0712 ( PRDP0712 ) ,.PRDP0709 ( PRDP0709 )
     ,.PRDP0708 ( PRDP0708 ) ,.PRDSCN15 ( PRDSCN15 ) ,.PRDSCN14 ( PRDSCN14 )
     ,.PRDSCN13 ( PRDSCN13 ) ,.PRDSCN12 ( PRDSCN12 ) ,.PSELCIB4 ( PSELCIB4 )
     ,.PRDSCN11 ( PRDSCN11 ) ,.PRDSCN10 ( PRDSCN10 ) ,.PSELFCB2 ( PSELFCB2 )
     ,.PRDSCN9 ( PRDSCN9 ) ,.PRDSCN8 ( PRDSCN8 ) ,.PRDSCN7 ( PRDSCN7 )
     ,.PRDSCN6 ( PRDSCN6 ) ,.PRDSCN5 ( PRDSCN5 ) ,.PRDSCN4 ( PRDSCN4 )
     ,.PRDSCN3 ( PRDSCN3 ) ,.PRDSCN2 ( PRDSCN2 ) ,.PRDSCN1 ( PRDSCN1 )
     ,.PRDSCN0 ( PRDSCN0 ) ,.PRDMAW15 ( PRDMAW15 ) ,.PRDMAW14 ( PRDMAW14 )
     ,.PRDMAW13 ( PRDMAW13 ) ,.PRDMAW12 ( PRDMAW12 ) ,.PRDMAW11 ( PRDMAW11 )
     ,.PRDMAW10 ( PRDMAW10 ) ,.PRDMAW9 ( PRDMAW9 ) ,.PRDMAW8 ( PRDMAW8 )
     ,.PRDMAW7 ( PRDMAW7 ) ,.PRDMAW6 ( PRDMAW6 ) ,.PRDMAW5 ( PRDMAW5 )
     ,.PRDMAW4 ( PRDMAW4 ) ,.PSELAD2 ( PSELAD2 ) ,.PRDMAW3 ( PRDMAW3 )
     ,.PSELAD1 ( PSELAD1 ) ,.PRDMAW2 ( PRDMAW2 ) ,.PRDMAW1 ( PRDMAW1 )
     ,.PRDMAW0 ( PRDMAW0 ) ,.PRDCRC15 ( PRDCRC15 ) ,.PRDCRC14 ( PRDCRC14 )
     ,.PRDCRC13 ( PRDCRC13 ) ,.PRDCRC12 ( PRDCRC12 ) ,.PRDCRC11 ( PRDCRC11 )
     ,.PRDCRC10 ( PRDCRC10 ) ,.PRDCRC3 ( PRDCRC3 ) ,.PRDCRC2 ( PRDCRC2 )
     ,.PRDCRC1 ( PRDCRC1 ) ,.PRDCRC0 ( PRDCRC0 ) ,.BBPRDATA15 ( BBPRDATA15 )
     ,.BBPRDATA14 ( BBPRDATA14 ) ,.BBPRDATA13 ( BBPRDATA13 ) ,.BBPRDATA12 ( BBPRDATA12 )
     ,.BBPRDATA11 ( BBPRDATA11 ) ,.BBPRDATA10 ( BBPRDATA10 ) ,.BBPRDATA9 ( BBPRDATA9 )
     ,.BBPRDATA8 ( BBPRDATA8 ) ,.BBPRDATA7 ( BBPRDATA7 ) ,.BBPRDATA6 ( BBPRDATA6 )
     ,.BBPRDATA5 ( BBPRDATA5 ) ,.BBPRDATA4 ( BBPRDATA4 ) ,.BBPRDATA3 ( BBPRDATA3 )
     ,.BBPRDATA2 ( BBPRDATA2 ) ,.BBPRDATA1 ( BBPRDATA1 ) ,.BBPRDATA0 ( BBPRDATA0 )
     ,.PWRITE ( PWRITE ) ,.BBPENABLE ( BBPENABLE ) ,.BBPWRITE ( BBPWRITE )
     ,.BBMA15 ( BBMA15 ) ,.BBMA14 ( BBMA14 ) ,.BBMA13 ( BBMA13 ) ,.BBMA12 ( BBMA12 )
     ,.BBMA11 ( BBMA11 ) ,.BBMA10 ( BBMA10 ) ,.BBMA9 ( BBMA9 ) ,.BBMA8 ( BBMA8 )
     ,.BBMA7 ( BBMA7 ) ,.BBMA6 ( BBMA6 ) ,.BBMA5 ( BBMA5 ) ,.BBMA4 ( BBMA4 )
     ,.BBMA3 ( BBMA3 ) ,.BBMA2 ( BBMA2 ) ,.BBMA1 ( BBMA1 ) ,.BBMA0 ( BBMA0 )
     ,.PADDR6 ( PADDR6 ) ,.PADDR5 ( PADDR5 ) ,.PADDR4 ( PADDR4 ) ,.PADDR3 ( PADDR3 )
     ,.PADDR2 ( PADDR2 ) ,.PADDR1 ( PADDR1 ) ,.PADDR0 ( PADDR0 ) ,.PSELP0 ( PSELP0 )
     ,.PSELP1 ( PSELP1 ) ,.PSELP2 ( PSELP2 ) ,.PSELP3 ( PSELP3 ) ,.PSELP4 ( PSELP4 )
     ,.PSELP5 ( PSELP5 ) ,.PSELP6 ( PSELP6 ) ,.PSELP7 ( PSELP7 ) ,.PSELP14 ( PSELP14 )
     ,.PSELSA01 ( PSELSA01 ) ,.PSELSA02 ( PSELSA02 ) ,.PSELSA11 ( PSELSA11 )
     ,.PSELSA12 ( PSELSA12 ) ,.PSELKR ( PSELKR ) ,.PSELIM8 ( PSELIM8 )
     ,.PSELIM4 ( PSELIM4 ) ,.PSELIIC1 ( PSELIIC1 ) ,.PSELIIC2 ( PSELIIC2 )
     ,.PSELTA01 ( PSELTA01 ) ,.PSELTA02 ( PSELTA02 ) ,.PSELOCD1 ( PSELOCD1 )
     ,.PSELRTC ( PSELRTC ) ,.PSELWWDT ( PSELWWDT ) ,.PSELPCL ( PSELPCL )
     ,.PSELCSC1 ( PSELCSC1 ) ,.PSELCSC2 ( PSELCSC2 ) ,.PSELCSC3 ( PSELCSC3 )
     ,.PSELCPU ( PSELCPU ) ,.PSELDMAC ( PSELDMAC ) ,.PSELINT1 ( PSELINT1 )
     ,.PSELMD1 ( PSELMD1 ) ,.PSELMD2 ( PSELMD2 ) ,.PSELMOD1 ( PSELMOD1 )
     ,.PSELMOD2 ( PSELMOD2 ) ,.PSELPOG1 ( PSELPOG1 ) ,.PSELPOG2 ( PSELPOG2 )
     ,.PSELSCN ( PSELSCN ) ,.PSELCRC ( PSELCRC ) ,.PSELFCB1 ( PSELFCB1 )
     ,.PSELCIBC ( PSELCIBC ) ,.PSELCIBD ( PSELCIBD ) ,.BBSELSFR1 ( BBSELSFR1 )
     ,.BBSELSFR2 ( BBSELSFR2 ) ,.SLAPB ( SLAPB ) ,.MDR15 ( MDR15 ) ,.MDR14 ( MDR14 )
     ,.MDR13 ( MDR13 ) ,.MDR12 ( MDR12 ) ,.MDR11 ( MDR11 ) ,.MDR10 ( MDR10 )
     ,.MDR9 ( MDR9 ) ,.MDR8 ( MDR8 ) ,.MDR7 ( MDR7 ) ,.MDR6 ( MDR6 ) ,.MDR5 ( MDR5 )
     ,.MDR4 ( MDR4 ) ,.MDR3 ( MDR3 ) ,.MDR2 ( MDR2 ) ,.MDR1 ( MDR1 ) ,.MDR0 ( MDR0 )
     ,.MDWFLRO15 ( MDWFLRO15 ) ,.MDWFLRO14 ( MDWFLRO14 ) ,.MDWFLRO13 ( MDWFLRO13 )
     ,.MDWFLRO12 ( MDWFLRO12 ) ,.MDWFLRO11 ( MDWFLRO11 ) ,.MDWFLRO10 ( MDWFLRO10 )
     ,.MDWFLRO9 ( MDWFLRO9 ) ,.MDWFLRO8 ( MDWFLRO8 ) ,.MDWFLRO7 ( MDWFLRO7 )
     ,.MDWFLRO6 ( MDWFLRO6 ) ,.MDWFLRO5 ( MDWFLRO5 ) ,.MDWFLRO4 ( MDWFLRO4 )
     ,.MDWFLRO3 ( MDWFLRO3 ) ,.MDWFLRO2 ( MDWFLRO2 ) ,.MDWFLRO1 ( MDWFLRO1 )
     ,.MDWFLRO0 ( MDWFLRO0 ) ,.GDPORT ( GDPORT ) ,.GDINT ( GDINT ) ,.GDCSC ( GDCSC )
    
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_2.0/_macro/_local/kx4_porga_mf3_v2.00/_library/100821/kx4_porga.hdl
  KX4_PORGA porga (
    .PCLKRW ( PCLKRW ) ,.RESB ( RESB ) ,.SYSRESB ( SYSRESB ) ,.TESTMOD ( TESTMOD )
     ,.PRDSELEN ( PRDSELEN ) ,.PSEL1 ( PSELPOG1 ) ,.PSEL2 ( PSELPOG2 )
     ,.MA3 ( MA3 ) ,.MA2 ( MA2 ) ,.MA1 ( MA1 ) ,.MA0 ( MA0 ) ,.CPUWR ( CPUWR )
     ,.CPURD ( CPURD ) ,.TIN05 ( TIN05 ) ,.R15KOUT ( R15KOUT ) ,.FSUB ( FSUB )
     ,.OSCOUTM ( OSCOUTM ) ,.TNFEN01 ( TNFEN01 ) ,.BBCLK ( BBCLKR ) ,.P137EXINA ( P137EXINA )
     ,.SIN10 ( SIN10 ) ,.TIN07 ( TIN07 ) ,.MDR15 ( MDRPOG15 ) ,.MDR14 ( MDRPOG14 )
     ,.MDR13 ( MDRPOG13 ) ,.MDR12 ( MDRPOG12 ) ,.IAWEN ( IAWEN ) ,.MDR11 ( MDRPOG11 )
     ,.MDR10 ( MDRPOG10 ) ,.MDR9 ( MDRPOG9 ) ,.MDR8 ( MDRPOG8 ) ,.MDR7 ( MDRPOG7 )
     ,.MDR6 ( MDRPOG6 ) ,.MDR5 ( MDRPOG5 ) ,.MDR4 ( MDRPOG4 ) ,.MDR3 ( MDRPOG3 )
     ,.MDR2 ( MDRPOG2 ) ,.MDR1 ( MDRPOG1 ) ,.MDR0 ( MDRPOG0 ) ,.STOPZ ( STOPZ )
     ,.CHMOD ( CHMOD ) ,.SNFEN20 ( SNFEN20 ) ,.SNFEN10 ( SNFEN10 ) ,.SNFEN00 ( SNFEN00 )
     ,.TNFEN07 ( TNFEN07 ) ,.TNFEN06 ( TNFEN06 ) ,.TNFEN05 ( TNFEN05 )
     ,.TNFEN04 ( TNFEN04 ) ,.TNFEN03 ( TNFEN03 ) ,.TNFEN02 ( TNFEN02 )
     ,.TNFEN00 ( TNFEN00 ) ,.PIOR7 ( PIOR7 ) ,.PIOR6 ( PIOR6 ) ,.PIOR5 ( PIOR5 )
     ,.PIOR4 ( PIOR4 ) ,.PIOR3 ( PIOR3 ) ,.PIOR2 ( PIOR2 ) ,.PIOR1 ( PIOR1 )
     ,.PIOR0 ( PIOR0 ) ,.GDRAM1 ( GDRAM1 ) ,.GDRAM0 ( GDRAM0 ) ,.GDPORT ( GDPORT )
     ,.GDINT ( GDINT ) ,.GDCSC ( GDCSC ) ,.TIN05O ( TIN05O ) ,.INTP0EG ( INTP0EG )
     ,.TIN07O ( TIN07O ) ,.SEL20P ( SEL20P ) ,.SEL24P ( SEL24P ) ,.SEL32P ( SEL32P )
     ,.SEL40P ( SEL40P ) ,.SEL08P ( SEL08P ) ,.SEL30P ( SEL30P ) ,.SEL36P ( SEL36P )
     ,.SEL44P ( SEL44P ) ,.SEL52P ( SEL52P ) ,.SEL38P ( SEL38P ) ,.SEL48P ( SEL48P )
     ,.SEL64P ( SEL64P ) ,.RAMSIZE7 ( RAMSIZE7ICE ) ,.RAMSIZE6 ( RAMSIZE6ICE )
     ,.RAMSIZE5 ( RAMSIZE5ICE ) ,.RAMSIZE4 ( RAMSIZE4ICE ) ,.RAMSIZE3 ( RAMSIZE3ICE )
     ,.RAMSIZE2 ( RAMSIZE2ICE ) ,.RAMSIZE1 ( RAMSIZE1ICE ) ,.RAMSIZE0 ( RAMSIZE0ICE )
     ,.FLSIZE3 ( FLSIZE3ICE ) ,.FLSIZE2 ( FLSIZE2ICE ) ,.FLSIZE1 ( FLSIZE1ICE )
     ,.FLSIZE0 ( FLSIZE0ICE ) ,.DFSIZE1 ( DFSIZE1ICE ) ,.DFSIZE0 ( DFSIZE0ICE )
     ,.SYSRSOUTB ( SYSRSOUTB ) ,.SEL20PI ( SEL20PI ) ,.SEL24PI ( SEL24PI )
     ,.SEL32PI ( SEL32PI ) ,.SEL40PI ( SEL40PI ) ,.SEL30PI ( SEL30PI )
     ,.SEL36PI ( SEL36PI ) ,.SEL44PI ( SEL44PI ) ,.SEL52PI ( SEL52PI )
     ,.SEL38PI ( SEL38PI ) ,.SEL48PI ( SEL48PI ) ,.SEL64PI ( SEL64PI )
     ,.MDWFLRO15 ( MDWFLRO15 ) ,.MDWFLRO14 ( MDWFLRO14 ) ,.MDWFLRO13 ( MDWFLRO13 )
     ,.MDWFLRO12 ( MDWFLRO12 ) ,.MDWFLRO11 ( MDWFLRO11 ) ,.MDWFLRO10 ( MDWFLRO10 )
     ,.MDWFLRO9 ( MDWFLRO9 ) ,.MDWFLRO8 ( MDWFLRO8 ) ,.MDWFLRO7 ( MDWFLRO7 )
     ,.MDWFLRO6 ( MDWFLRO6 ) ,.MDWFLRO5 ( MDWFLRO5 ) ,.MDWFLRO4 ( MDWFLRO4 )
     ,.MDWFLRO3 ( MDWFLRO3 ) ,.MDWFLRO2 ( MDWFLRO2 ) ,.MDWFLRO1 ( MDWFLRO1 )
     ,.MDWFLRO0 ( MDWFLRO0 ) ,.DGEN07 ( DGEN07 ) ,.DGEN06 ( DGEN06 ) ,.DGEN05 ( DGEN05 )
     ,.DGEN04 ( DGEN04 ) ,.DGEN03 ( DGEN03 ) ,.DGEN02 ( DGEN02 ) ,.DGEN01 ( DGEN01 )
     ,.DGEN00 ( DGEN00 ) ,.SCANMODE ( SCANMODE ) ,.BBISC ( BBISC ) ,.SIN00 ( SIN00 )
    
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_2.0/_macro/_local/kx4_intor_mf3_v2.00/_library/101207/kx4_intor.hdl
  KX4_INTOR intor (
    .INTSRE0 ( INTSRE0 ) ,.INTTM01H ( INTTM01H ) ,.INTSRE1 ( INTSRE1 )
     ,.INTTM03H ( INTTM03H ) ,.INTP6 ( INTP6 ) ,.INTP7 ( INTP7 ) ,.INTP8 ( INTP8 )
     ,.INTP9 ( INTP9 ) ,.INTP10 ( INTP10 ) ,.INTP11 ( INTP11 ) ,.BBINT3 ( BBINT3 )
     ,.BBINT4 ( BBINT4 ) ,.BBINT5 ( BBINT5 ) ,.BBINT6 ( BBINT6 ) ,.BBINT7 ( BBINT7 )
     ,.BBINT8 ( BBINT8 ) ,.INTAS22 ( INTAS22 ) ,.INTAS28 ( INTAS28 ) ,.INTAS52 ( INTAS52 )
     ,.INTAS4A ( INTAS4A ) ,.INTAS4C ( INTAS4C ) ,.INTAS4E ( INTAS4E )
     ,.INTAS50 ( INTAS50 ) ,.INTAS54 ( INTAS54 ) ,.INTWWDT ( INTWWDT )
     ,.INTSRO ( INTSRO ) ,.INTAS04 ( INTAS04 )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_1.0/_macro/_local/kx4_ckdist_mf3_v1.00/_library/100130/kx4_ckdist.hdl
  KX4_CKDIST ckdist (
    .PRSCLK1 ( PRSCLK1 ) ,.PRSCLK2 ( PRSCLK2 ) ,.PRSCLK3 ( PRSCLK3 ) ,.PRSCLK4 ( PRSCLK4 )
     ,.PRSCLK5 ( PRSCLK5 ) ,.PRSCLK6 ( PRSCLK6 ) ,.PRSCLK7 ( PRSCLK7 )
     ,.PRSCLK8 ( PRSCLK8 ) ,.PRSCLK9 ( PRSCLK9 ) ,.PRSCLK10 ( PRSCLK10 )
     ,.PRSCLK11 ( PRSCLK11 ) ,.PRSCLK12 ( PRSCLK12 ) ,.PRSCLK13 ( PRSCLK13 )
     ,.PRSCLK14 ( PRSCLK14 ) ,.PRSCLK15 ( PRSCLK15 ) ,.PRST003 ( PRST003 )
     ,.PRST011 ( PRST011 ) ,.PRST002 ( PRST002 ) ,.PRST010 ( PRST010 )
     ,.PRST001 ( PRST001 ) ,.PRSS113 ( PRSS113 ) ,.PRST000 ( PRST000 )
     ,.PRSS112 ( PRSS112 ) ,.PRST013 ( PRST013 ) ,.PRST021 ( PRST021 )
     ,.PRST012 ( PRST012 ) ,.PRST020 ( PRST020 ) ,.PRST031 ( PRST031 )
     ,.PRST030 ( PRST030 ) ,.PRSS003 ( PRSS003 ) ,.PRSS011 ( PRSS011 )
     ,.PRSS002 ( PRSS002 ) ,.PRSS010 ( PRSS010 ) ,.PRSS001 ( PRSS001 )
     ,.PRSS000 ( PRSS000 ) ,.PRSS013 ( PRSS013 ) ,.PRSS101 ( PRSS101 )
     ,.PRSS012 ( PRSS012 ) ,.PRSS100 ( PRSS100 ) ,.PRSS103 ( PRSS103 )
     ,.PRSS111 ( PRSS111 ) ,.PRSS102 ( PRSS102 ) ,.PRSS110 ( PRSS110 )
     ,.PRSI000 ( PRSI000 ) ,.CK0TAU0 ( CK0TAU0 ) ,.CK1TAU0 ( CK1TAU0 )
     ,.CK2TAU0 ( CK2TAU0 ) ,.CK3TAU0 ( CK3TAU0 ) ,.CK0SAU0 ( CK0SAU0 )
     ,.CK1SAU0 ( CK1SAU0 ) ,.CK0SAU1 ( CK0SAU1 ) ,.CK1SAU1 ( CK1SAU1 )
     ,.CK0IIC0 ( CK0IIC0 ) ,.SVPERI0 ( SVPERI0 ) ,.SVPERI1 ( SVPERI1 )
    
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_1.0/_macro/_local/kx4_monsig_mf3_v1.00/_library/100202/kx4_monsig.hdl
  KX4_MONSIG monsig (
    .R32MOUT ( R32MOUT ) ,.R15KOUT ( R15KOUT ) ,.FIHFL ( FIHFL ) ,.FIHOCD ( FIHOCD )
     ,.TR32MOUT ( TR32MOUT ) ,.TR15KOUT ( TR15KOUT ) ,.TFIHFL ( TFIHFL )
     ,.TFIHOCD ( TFIHOCD ) ,.TESTMOD ( TESTMOD )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_1.0/_macro/_soft/qlk0rintm4v1_mf3_v1.00/_library/_df3.0_100206/qlk0rintm4v1.hdl_100206
  QLK0RINTM4V1 intm4 (
    .MDR11 ( MDRIM411 ) ,.MDR10 ( MDRIM410 ) ,.MDR9 ( MDRIM49 ) ,.MDR8 ( MDRIM48 )
     ,.MDR3 ( MDRIM43 ) ,.MDR2 ( MDRIM42 ) ,.MDR1 ( MDRIM41 ) ,.MDR0 ( MDRIM40 )
     ,.MDW11 ( MDW11 ) ,.MDW10 ( MDW10 ) ,.MDW9 ( MDW9 ) ,.MDW8 ( MDW8 )
     ,.MDW3 ( MDW3 ) ,.MDW2 ( MDW2 ) ,.MDW1 ( MDW1 ) ,.MDW0 ( MDW0 ) ,.MA0 ( MA0 )
     ,.PCLKRW ( PCLKRW ) ,.PSELINTM ( PSELIM4 ) ,.CPURD ( CPURD ) ,.CPUWR ( CPUWR )
     ,.RESB ( RESB ) ,.INTP3 ( INTP11 ) ,.INTP2 ( INTP10 ) ,.INTP1 ( INTP9 )
     ,.INTP0 ( INTP8 ) ,.EGIN3 ( INTP11EG ) ,.EGIN2 ( INTP10EG ) ,.EGIN1 ( P75EXINA )
     ,.EGIN0 ( P74EXINA ) ,.SVMOD ( SVPERI1 ) ,.SCANMODE ( SCANMODE ) ,.ICECK60M ( ICECK60M )
    
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_1.0/_macro/_soft/qlk0rintm8v1_mf3_v1.00/_library/_df3.0_100206/qlk0rintm8v1.hdl_100206
  QLK0RINTM8V1 intm8 (
    .MDR15 ( MDRIM815 ) ,.MDR14 ( MDRIM814 ) ,.MDR13 ( MDRIM813 ) ,.MDR12 ( MDRIM812 )
     ,.MDR11 ( MDRIM811 ) ,.MDR10 ( MDRIM810 ) ,.MDR9 ( MDRIM89 ) ,.MDR8 ( MDRIM88 )
     ,.MDR7 ( MDRIM87 ) ,.MDR6 ( MDRIM86 ) ,.MDR5 ( MDRIM85 ) ,.MDR4 ( MDRIM84 )
     ,.MDR3 ( MDRIM83 ) ,.MDR2 ( MDRIM82 ) ,.MDR1 ( MDRIM81 ) ,.MDR0 ( MDRIM80 )
     ,.MDW15 ( MDW15 ) ,.MDW14 ( MDW14 ) ,.MDW13 ( MDW13 ) ,.MDW12 ( MDW12 )
     ,.MDW11 ( MDW11 ) ,.MDW10 ( MDW10 ) ,.MDW9 ( MDW9 ) ,.MDW8 ( MDW8 )
     ,.MDW7 ( MDW7 ) ,.MDW6 ( MDW6 ) ,.MDW5 ( MDW5 ) ,.MDW4 ( MDW4 ) ,.MDW3 ( MDW3 )
     ,.MDW2 ( MDW2 ) ,.MDW1 ( MDW1 ) ,.MDW0 ( MDW0 ) ,.MA0 ( MA0 ) ,.PCLKRW ( PCLKRW )
     ,.PSELINTM ( PSELIM8 ) ,.CPURD ( CPURD ) ,.CPUWR ( CPUWR ) ,.RESB ( RESB )
     ,.INTP7 ( INTP7 ) ,.INTP6 ( INTP6 ) ,.INTP5 ( INTP5 ) ,.INTP4 ( INTP4 )
     ,.INTP3 ( INTP3 ) ,.INTP2 ( INTP2 ) ,.INTP1 ( INTP1 ) ,.INTP0 ( INTP0 )
     ,.EGIN7 ( P141EXINA ) ,.EGIN6 ( P140EXINA ) ,.EGIN5 ( INTP5EG ) ,.EGIN4 ( P31EXINA )
     ,.EGIN3 ( P30EXINA ) ,.EGIN2 ( P51EXINA ) ,.EGIN1 ( P50EXINA ) ,.EGIN0 ( INTP0EG )
     ,.SVMOD ( SVPERI1 ) ,.SCANMODE ( SCANMODE ) ,.ICECK60M ( ICECK60M )
    
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_2.0/_macro/_local/kx4_iicascldly_mf3_v1.10/_library/101105/kx4_iicascldly.hdl
  KX4_IICASCLDLY sdadly0 (
    .SCL ( SCLI0 ) ,.SCLDLY ( SCLI1DLY ) ,.SCANMODE ( SCANMODE ) ,.CLK60M ( CLK60M )
    
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/_ice/_macro/_zantei/_iicasdadly_20101111/kx4_iicasdadly.hdl
  KX4_IICASDADLY sdadly1 (
    .SDA ( SDAI0 ) ,.SDADLY ( SDAI1DLY ) ,.SCANMODE ( SCANMODE ) ,.CLK60M ( CLK60M )
    
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_1.0/_macro/_local/kx4_sdadly_mf3_v1.00/_library/100218/kx4_sdadly.hdl
  KX4_SDADLY sdadly2 (
    .SOUT ( SOUT012 ) ,.SOUTDLY ( SOUT012DLY ) ,.SCANMODE ( SCANMODE )
     ,.CLK60M ( CLK60M )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_1.0/_macro/_local/kx4_sdadly_mf3_v1.00/_library/100218/kx4_sdadly.hdl
  KX4_SDADLY sdadly3 (
    .SOUT ( SOUT010 ) ,.SOUTDLY ( SOUT010DLY ) ,.SCANMODE ( SCANMODE )
     ,.CLK60M ( CLK60M )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_1.0/_macro/_local/kx4_sdadly_mf3_v1.00/_library/100218/kx4_sdadly.hdl
  KX4_SDADLY sdadly011 (
    .SOUT ( SOUT011 ) ,.SOUTDLY ( SOUT011DLY ) ,.SCANMODE ( SCANMODE )
     ,.CLK60M ( CLK60M )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_1.0/_macro/_local/kx4_sdadly_mf3_v1.00/_library/100218/kx4_sdadly.hdl
  KX4_SDADLY sdadly013 (
    .SOUT ( SOUT013 ) ,.SOUTDLY ( SOUT013DLY ) ,.SCANMODE ( SCANMODE )
     ,.CLK60M ( CLK60M )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_1.0/_macro/_local/kx4_sdadly_mf3_v1.00/_library/100218/kx4_sdadly.hdl
  KX4_SDADLY sdadly110 (
    .SOUT ( SOUT110 ) ,.SOUTDLY ( SOUT110DLY ) ,.SCANMODE ( SCANMODE )
     ,.CLK60M ( CLK60M )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_1.0/_macro/_local/kx4_sdadly_mf3_v1.00/_library/100218/kx4_sdadly.hdl
  KX4_SDADLY sdadly111 (
    .SOUT ( SOUT111 ) ,.SOUTDLY ( SOUT111DLY ) ,.SCANMODE ( SCANMODE )
     ,.CLK60M ( CLK60M )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_1.0/_macro/_soft/qlk0riicav2_mf3_v2.00/_library/QLK0RIICAV2.v
  QLK0RIICAV2 iica (
    .PCLK ( PCLKIIC ) ,.PCLKRW ( PCLKRW ) ,.PRESETZ ( PRESIICZ ) ,.CK0 ( CK0IIC0 )
     ,.SCANCLK ( SCANCLK ) ,.PADDR2 ( PADDR2 ) ,.PADDR1 ( PADDR1 ) ,.PADDR0 ( PADDR0 )
     ,.PWDATA15 ( MDW15 ) ,.PWDATA14 ( MDW14 ) ,.PWDATA13 ( MDW13 ) ,.PWDATA12 ( MDW12 )
     ,.PWDATA11 ( MDW11 ) ,.PWDATA10 ( MDW10 ) ,.PWDATA9 ( MDW9 ) ,.PWDATA8 ( MDW8 )
     ,.PWDATA7 ( MDW7 ) ,.PWDATA6 ( MDW6 ) ,.PWDATA5 ( MDW5 ) ,.PWDATA4 ( MDW4 )
     ,.PWDATA3 ( MDW3 ) ,.PWDATA2 ( MDW2 ) ,.PWDATA1 ( MDW1 ) ,.PWDATA0 ( MDW0 )
     ,.PRDATA15 ( PRDIIC15 ) ,.PRDATA14 ( PRDIIC14 ) ,.PRDATA13 ( PRDIIC13 )
     ,.PRDATA12 ( PRDIIC12 ) ,.PRDATA11 ( PRDIIC11 ) ,.PRDATA10 ( PRDIIC10 )
     ,.PRDATA9 ( PRDIIC9 ) ,.PRDATA8 ( PRDIIC8 ) ,.PRDATA7 ( PRDIIC7 )
     ,.PRDATA6 ( PRDIIC6 ) ,.PRDATA5 ( PRDIIC5 ) ,.PRDATA4 ( PRDIIC4 )
     ,.PRDATA3 ( PRDIIC3 ) ,.PRDATA2 ( PRDIIC2 ) ,.PRDATA1 ( PRDIIC1 )
     ,.PRDATA0 ( PRDIIC0 ) ,.PWRITE ( PWRITE ) ,.PENABLE ( PENABLE ) ,.PSEL1 ( PSELIIC2 )
     ,.PSEL0 ( PSELIIC1 ) ,.SCANMODE ( SCANMODE ) ,.SVMOD ( SVPERI1 ) ,.PRS0 ( PRSI000 )
     ,.SCLI0 ( SCLI0 ) ,.SCLI1 ( SCLI1DLY ) ,.SDAI0 ( SDAI0 ) ,.SDAI1 ( SDAI1DLY )
     ,.SCLO0 ( SCLO0 ) ,.SDAO0 ( SDAO0 ) ,.SCLO1 ( SCLO1 ) ,.SDAO1 ( SDAO1 )
     ,.INTIIC0 ( INTIIC0 ) ,.SCANEN ( SCANEN )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_1.0/_macro/_soft/qlk0rsau04r2v1_mf3_v1.00/_library/QLK0RSAU04R2V1.v
  QLK0RSAU04R2V1 sau0 (
    .PCLK ( PCLKSAU0 ) ,.PCLKRW ( PCLKRW ) ,.PRESETZ ( PRESSAU0Z ) ,.PSEL2 ( PSELSA02 )
     ,.PSEL1 ( PSELSA01 ) ,.PENABLE ( PENABLE ) ,.PWRITE ( PWRITE ) ,.PADDR5 ( PADDR5 )
     ,.PADDR4 ( PADDR4 ) ,.PADDR3 ( PADDR3 ) ,.PADDR2 ( PADDR2 ) ,.PADDR1 ( PADDR1 )
     ,.PWDATA31 ( MDW15 ) ,.PWDATA23 ( MDW7 ) ,.PWDATA15 ( MDW15 ) ,.PWDATA30 ( MDW14 )
     ,.PWDATA22 ( MDW6 ) ,.PWDATA14 ( MDW14 ) ,.PWDATA29 ( MDW13 ) ,.PWDATA28 ( MDW12 )
     ,.PWDATA27 ( MDW11 ) ,.PWDATA19 ( MDW3 ) ,.PWDATA26 ( MDW10 ) ,.PWDATA18 ( MDW2 )
     ,.PWDATA25 ( MDW9 ) ,.PWDATA17 ( MDW1 ) ,.PWDATA24 ( MDW8 ) ,.PWDATA16 ( MDW0 )
     ,.PWDATA21 ( MDW5 ) ,.PWDATA13 ( MDW13 ) ,.PWDATA20 ( MDW4 ) ,.PWDATA12 ( MDW12 )
     ,.PWDATA11 ( MDW11 ) ,.PWDATA10 ( MDW10 ) ,.PWDATA9 ( MDW9 ) ,.PWDATA8 ( MDW8 )
     ,.PWDATA7 ( MDW7 ) ,.PWDATA6 ( MDW6 ) ,.PWDATA5 ( MDW5 ) ,.PWDATA4 ( MDW4 )
     ,.PWDATA3 ( MDW3 ) ,.PWDATA2 ( MDW2 ) ,.PWDATA1 ( MDW1 ) ,.PWDATA0 ( MDW0 )
     ,.PRDATA15 ( PRDSA015 ) ,.PRDATA14 ( PRDSA014 ) ,.PRDATA13 ( PRDSA013 )
     ,.PRDATA12 ( PRDSA012 ) ,.PRDATA11 ( PRDSA011 ) ,.PRDATA10 ( PRDSA010 )
     ,.PRDATA9 ( PRDSA09 ) ,.PRDATA8 ( PRDSA08 ) ,.PRDATA7 ( PRDSA07 )
     ,.PRDATA6 ( PRDSA06 ) ,.PRDATA5 ( PRDSA05 ) ,.PRDATA4 ( PRDSA04 )
     ,.PRDATA3 ( PRDSA03 ) ,.PRDATA2 ( PRDSA02 ) ,.PRDATA1 ( PRDSA01 )
     ,.PRDATA0 ( PRDSA00 ) ,.INT0 ( INTSAU00 ) ,.INT1 ( INTSAU01 ) ,.SEINT0 ( SEINT0SAU0 )
     ,.SEINT1 ( INTSRE0 ) ,.SIN0 ( SIN00 ) ,.SIN1 ( P74EXINA ) ,.SOUT00 ( SOUT000 )
     ,.SOUT01 ( SOUT001 ) ,.SOUT10 ( SOUT010 ) ,.SOUT02 ( SOUT002 ) ,.SOUT11 ( SOUT011 )
     ,.SOUT03 ( SOUT003 ) ,.SCKO0 ( SCKO00 ) ,.SCKO1 ( SCKO01 ) ,.SCKI0 ( SCKI00 )
     ,.SCKI1 ( P75EXINA ) ,.NFEN0 ( SNFEN00 ) ,.INT2 ( INTSAU02 ) ,.INT3 ( INTSAU03 )
     ,.SEINT2 ( SEINT2SAU0 ) ,.SEINT3 ( INTSRE1 ) ,.SIN2 ( SIN02 ) ,.SIN3 ( SIN03 )
     ,.SOUT12 ( SOUT012 ) ,.SOUT13 ( SOUT013 ) ,.SCKO2 ( SCKO02 ) ,.SCKO3 ( SCKO03 )
     ,.SCKI2 ( P04EXINA ) ,.SCKI3 ( P30EXINA ) ,.NFEN2 ( SNFEN10 ) ,.PRS13 ( PRSS013 )
     ,.PRS12 ( PRSS012 ) ,.PRS11 ( PRSS011 ) ,.PRS03 ( PRSS003 ) ,.PRS10 ( PRSS010 )
     ,.PRS02 ( PRSS002 ) ,.PRS01 ( PRSS001 ) ,.PRS00 ( PRSS000 ) ,.CK0 ( CK0SAU0 )
     ,.CK1 ( CK1SAU0 ) ,.REQPCLK ( REQPCLKSAU0 ) ,.SCANEN ( SCANEN ) ,.SCANMODE ( SCANMODE )
    
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_1.0/_macro/_soft/qlk0rsau02r2v1_mf3_v1.00/_library/QLK0RSAU02R2V1.v
  QLK0RSAU02R2V1 sau1 (
    .PCLK ( PCLKSAU1 ) ,.PCLKRW ( PCLKRW ) ,.PRESETZ ( PRESSAU1Z ) ,.PSEL2 ( PSELSA12 )
     ,.PSEL1 ( PSELSA11 ) ,.PENABLE ( PENABLE ) ,.PWRITE ( PWRITE ) ,.PADDR5 ( PADDR5 )
     ,.PADDR4 ( PADDR4 ) ,.PADDR3 ( PADDR3 ) ,.PADDR2 ( PADDR2 ) ,.PADDR1 ( PADDR1 )
     ,.PWDATA31 ( MDW15 ) ,.PWDATA23 ( MDW7 ) ,.PWDATA15 ( MDW15 ) ,.PWDATA30 ( MDW14 )
     ,.PWDATA22 ( MDW6 ) ,.PWDATA14 ( MDW14 ) ,.PWDATA29 ( MDW13 ) ,.PWDATA28 ( MDW12 )
     ,.PWDATA27 ( MDW11 ) ,.PWDATA19 ( MDW3 ) ,.PWDATA26 ( MDW10 ) ,.PWDATA18 ( MDW2 )
     ,.PWDATA25 ( MDW9 ) ,.PWDATA17 ( MDW1 ) ,.PWDATA24 ( MDW8 ) ,.PWDATA16 ( MDW0 )
     ,.PWDATA21 ( MDW5 ) ,.PWDATA13 ( MDW13 ) ,.PWDATA20 ( MDW4 ) ,.PWDATA12 ( MDW12 )
     ,.PWDATA11 ( MDW11 ) ,.PWDATA10 ( MDW10 ) ,.PWDATA9 ( MDW9 ) ,.PWDATA8 ( MDW8 )
     ,.PWDATA7 ( MDW7 ) ,.PWDATA6 ( MDW6 ) ,.PWDATA5 ( MDW5 ) ,.PWDATA4 ( MDW4 )
     ,.PWDATA3 ( MDW3 ) ,.PWDATA2 ( MDW2 ) ,.PWDATA1 ( MDW1 ) ,.PWDATA0 ( MDW0 )
     ,.PRDATA15 ( PRDSA115 ) ,.PRDATA14 ( PRDSA114 ) ,.PRDATA13 ( PRDSA113 )
     ,.PRDATA12 ( PRDSA112 ) ,.PRDATA11 ( PRDSA111 ) ,.PRDATA10 ( PRDSA110 )
     ,.PRDATA9 ( PRDSA19 ) ,.PRDATA8 ( PRDSA18 ) ,.PRDATA7 ( PRDSA17 )
     ,.PRDATA6 ( PRDSA16 ) ,.PRDATA5 ( PRDSA15 ) ,.PRDATA4 ( PRDSA14 )
     ,.PRDATA3 ( PRDSA13 ) ,.PRDATA2 ( PRDSA12 ) ,.PRDATA1 ( PRDSA11 )
     ,.PRDATA0 ( PRDSA10 ) ,.INT0 ( INTSAU10 ) ,.INT1 ( INTSAU11 ) ,.SEINT0 ( SEINT0SAU1 )
     ,.SEINT1 ( INTSRE2 ) ,.SIN0 ( SIN10 ) ,.SIN1 ( P71EXINA ) ,.SOUT00 ( SOUT100 )
     ,.SOUT01 ( SOUT101 ) ,.SOUT10 ( SOUT110 ) ,.SOUT11 ( SOUT111 ) ,.SCKO0 ( SCKO10 )
     ,.SCKO1 ( SCKO11 ) ,.SCKI0 ( P15EXINA ) ,.SCKI1 ( P70EXINA ) ,.NFEN0 ( SNFEN20 )
     ,.PRS13 ( PRSS113 ) ,.PRS12 ( PRSS112 ) ,.PRS11 ( PRSS111 ) ,.PRS03 ( PRSS103 )
     ,.PRS10 ( PRSS110 ) ,.PRS02 ( PRSS102 ) ,.PRS01 ( PRSS101 ) ,.PRS00 ( PRSS100 )
     ,.CK0 ( CK0SAU1 ) ,.CK1 ( CK1SAU1 ) ,.SCANEN ( SCANEN ) ,.SCANMODE ( SCANMODE )
    
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_1.0/_macro/_soft/qlk0rtau08r2v1_mf3_v1.00/_library/QLK0RTAU08R2V1.v
  QLK0RTAU08R2V1 tau0 (
    .PCLK ( PCLKTAU0 ) ,.PCLKRW ( PCLKRW ) ,.PRESETZ ( PRESTAU0Z ) ,.PSEL2 ( PSELTA02 )
     ,.PSEL1 ( PSELTA01 ) ,.PADDR5 ( PADDR5 ) ,.PADDR4 ( PADDR4 ) ,.PADDR3 ( PADDR3 )
     ,.PADDR2 ( PADDR2 ) ,.PADDR1 ( PADDR1 ) ,.PADDR0 ( PADDR0 ) ,.PENABLE ( PENABLE )
     ,.PWRITE ( PWRITE ) ,.PWDATA31 ( MDW15 ) ,.PWDATA23 ( MDW7 ) ,.PWDATA15 ( MDW15 )
     ,.PWDATA30 ( MDW14 ) ,.PWDATA22 ( MDW6 ) ,.PWDATA14 ( MDW14 ) ,.PWDATA29 ( MDW13 )
     ,.PWDATA28 ( MDW12 ) ,.PWDATA27 ( MDW11 ) ,.PWDATA19 ( MDW3 ) ,.PWDATA26 ( MDW10 )
     ,.PWDATA18 ( MDW2 ) ,.PWDATA25 ( MDW9 ) ,.PWDATA17 ( MDW1 ) ,.PWDATA24 ( MDW8 )
     ,.PWDATA16 ( MDW0 ) ,.PWDATA21 ( MDW5 ) ,.PWDATA13 ( MDW13 ) ,.PWDATA20 ( MDW4 )
     ,.PWDATA12 ( MDW12 ) ,.PWDATA11 ( MDW11 ) ,.PWDATA10 ( MDW10 ) ,.PWDATA9 ( MDW9 )
     ,.PWDATA8 ( MDW8 ) ,.PWDATA7 ( MDW7 ) ,.PWDATA6 ( MDW6 ) ,.PWDATA5 ( MDW5 )
     ,.PWDATA4 ( MDW4 ) ,.PWDATA3 ( MDW3 ) ,.PWDATA2 ( MDW2 ) ,.PWDATA1 ( MDW1 )
     ,.PWDATA0 ( MDW0 ) ,.PRDATA15 ( PRDTA015 ) ,.PRDATA14 ( PRDTA014 )
     ,.PRDATA13 ( PRDTA013 ) ,.PRDATA12 ( PRDTA012 ) ,.PRDATA11 ( PRDTA011 )
     ,.PRDATA10 ( PRDTA010 ) ,.PRDATA9 ( PRDTA09 ) ,.PRDATA8 ( PRDTA08 )
     ,.PRDATA7 ( PRDTA07 ) ,.PRDATA6 ( PRDTA06 ) ,.PRDATA5 ( PRDTA05 )
     ,.PRDATA4 ( PRDTA04 ) ,.PRDATA3 ( PRDTA03 ) ,.PRDATA2 ( PRDTA02 )
     ,.PRDATA1 ( PRDTA01 ) ,.PRDATA0 ( PRDTA00 ) ,.CK3 ( CK3TAU0 ) ,.CK2 ( CK2TAU0 )
     ,.CK1 ( CK1TAU0 ) ,.CK0 ( CK0TAU0 ) ,.TIN7 ( TIN07O ) ,.TOE1 ( TOE01 )
     ,.TIN6 ( TIN06 ) ,.TOE0 ( TOE00 ) ,.TIN5 ( TIN05O ) ,.TIN4 ( TIN04 )
     ,.TIN3 ( TIN03 ) ,.TIN2 ( TIN02 ) ,.TIN1 ( P16EXINA ) ,.TIN0 ( OTI00 )
     ,.NFEN7 ( TNFEN07 ) ,.NFEN6 ( TNFEN06 ) ,.NFEN5 ( TNFEN05 ) ,.NFEN4 ( TNFEN04 )
     ,.NFEN3 ( TNFEN03 ) ,.NFEN2 ( TNFEN02 ) ,.NFEN1 ( TNFEN01 ) ,.NFEN0 ( TNFEN00 )
     ,.TOUT7 ( TOUT07 ) ,.TOUT6 ( TOUT06 ) ,.TOUT5 ( TOUT05 ) ,.TOUT4 ( TOUT04 )
     ,.TOUT3 ( TOUT03 ) ,.TOUT2 ( TOUT02 ) ,.TOUT1 ( TOUT01 ) ,.TOUT0 ( TOUT00 )
     ,.INT7 ( INTTM07 ) ,.INT6 ( INTTM06 ) ,.INT5 ( INTTM05 ) ,.INT4 ( INTTM04 )
     ,.INT3 ( INTTM03 ) ,.INT2 ( INTTM02 ) ,.INT1 ( INTTM01 ) ,.INT0 ( INTTM00 )
     ,.INTH3 ( INTTM03H ) ,.INTH1 ( INTTM01H ) ,.PRS31 ( PRST031 ) ,.PRS30 ( PRST030 )
     ,.PRS21 ( PRST021 ) ,.PRS13 ( PRST013 ) ,.PRS20 ( PRST020 ) ,.PRS12 ( PRST012 )
     ,.PRS11 ( PRST011 ) ,.PRS03 ( PRST003 ) ,.PRS10 ( PRST010 ) ,.PRS02 ( PRST002 )
     ,.PRS01 ( PRST001 ) ,.PRS00 ( PRST000 ) ,.CKEN7 ( CKENTAU07 ) ,.CKEN6 ( CKENTAU06 )
     ,.CKEN5 ( CKENTAU05 ) ,.CKEN4 ( CKENTAU04 ) ,.CKEN3 ( CKENTAU03 )
     ,.CKEN2 ( CKENTAU02 ) ,.CKEN1 ( CKENTAU01 ) ,.CKEN0 ( CKENTAU00 )
     ,.CDEN7 ( CDEN7 ) ,.CDEN6 ( CDEN6 ) ,.CDEN5 ( CDEN5 ) ,.CDEN4 ( CDEN4 )
     ,.CDEN3 ( CDEN3 ) ,.CDEN2 ( CDEN2 ) ,.CDEN1 ( CDEN1 ) ,.CDEN0 ( CDEN0 )
     ,.TOE7 ( TOE07 ) ,.TOE6 ( TOE06 ) ,.TOE5 ( TOE05 ) ,.TOE4 ( TOE04 )
     ,.TOE3 ( TOE03 ) ,.TOE2 ( TOE02 ) ,.TE7 ( TE07 ) ,.TE6 ( TE06 ) ,.TE5 ( TE05 )
     ,.TE4 ( TE04 ) ,.TE3 ( TE03 ) ,.TE2 ( TE02 ) ,.TE1 ( TE01 ) ,.TE0 ( TE00 )
    
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_2.0/_macro/_local/kx4_port0v1_mf3_v1.10/_library/100701/kx4_port0v1.hdl
  KX4_PORT0V1 port0 (
    .PCLKRW ( PCLKRW ) ,.PRESETZ ( RESB ) ,.PSEL ( PSELP0 ) ,.PWRITE ( PWRITE )
     ,.PENABLE ( PENABLE ) ,.PADDR4 ( PADDR4 ) ,.PADDR5 ( PADDR5 ) ,.PADDR6 ( PADDR6 )
     ,.PWDATA0 ( MDW0 ) ,.PWDATA1 ( MDW1 ) ,.PWDATA2 ( MDW2 ) ,.PWDATA3 ( MDW3 )
     ,.PWDATA4 ( MDW4 ) ,.PWDATA5 ( MDW5 ) ,.PWDATA6 ( MDW6 ) ,.NSRESB ( NSRESB )
     ,.SEL64P ( SEL64P ) ,.SEL48P ( SEL48P ) ,.SEL52P ( SEL52P ) ,.SEL44P ( SEL44P )
     ,.SEL36P ( SEL36P ) ,.SEL40P ( SEL40P ) ,.SEL32P ( SEL32P ) ,.SEL24P ( SEL24P )
     ,.SEL08P ( SEL08P ) ,.SEL38P ( SEL38P ) ,.SEL30P ( SEL30P ) ,.SEL20P ( SEL20P )
     ,.SEL64PI ( SEL64PI ) ,.SEL48PI ( SEL48PI ) ,.SEL52PI ( SEL52PI )
     ,.SEL44PI ( SEL44PI ) ,.SEL36PI ( SEL36PI ) ,.SEL40PI ( SEL40PI )
     ,.SEL32PI ( SEL32PI ) ,.SEL24PI ( SEL24PI ) ,.SEL38PI ( SEL38PI )
     ,.SEL30PI ( SEL30PI ) ,.SEL20PI ( SEL20PI ) ,.SCANMODE ( SCANMODE )
     ,.SCANCLK ( SCANCLK ) ,.TESDBT ( TESDBT2 ) ,.OPTOPLRD ( OPTOPLRD )
     ,.PRDATA0 ( PRDP0000 ) ,.PRDATA1 ( PRDP0001 ) ,.PRDATA2 ( PRDP0002 )
     ,.PRDATA3 ( PRDP0003 ) ,.PRDATA4 ( PRDP0004 ) ,.PRDATA5 ( PRDP0005 )
     ,.PRDATA6 ( PRDP0006 ) ,.PRDATA7 ( PRDP0007 ) ,.EXINA0 ( P00EXINA )
     ,.EXINA1 ( P01EXINA ) ,.EXINA2 ( P02EXINA ) ,.EXINA3 ( P03EXINA )
     ,.EXINA4 ( P04EXINA ) ,.EXINA5 ( P05EXINA ) ,.EXINA6 ( P06EXINA )
     ,.EXOUTA0 ( P00EXOUTA ) ,.EXOUTA1 ( pull_up60 ) ,.EXOUTA2 ( P02EXOUTA )
     ,.EXOUTB0 ( pull_down62 ) ,.EXOUTA3 ( SOUT012DLY ) ,.EXOUTB1 ( P01EXOUTB )
     ,.EXOUTA4 ( SCKO02 ) ,.EXOUTB2 ( pull_down65 ) ,.EXOUTC0 ( pull_down63 )
     ,.EXOUTA5 ( pull_up61 ) ,.EXOUTB3 ( P03EXOUTB ) ,.EXOUTC1 ( pull_down64 )
     ,.EXOUTA6 ( pull_up62 ) ,.EXOUTB4 ( pull_down68 ) ,.EXOUTC2 ( pull_down66 )
     ,.EXOUTB5 ( P05EXOUTB ) ,.EXOUTC3 ( pull_down67 ) ,.EXOUTB6 ( P06EXOUTB )
     ,.EXOUTC4 ( pull_down69 ) ,.EXOUTC5 ( pull_down70 ) ,.EXOUTC6 ( pull_down71 )
     ,.P00DIN ( P00DIN ) ,.P01DIN ( P01DIN ) ,.P02DIN ( P02DIN ) ,.P03DIN ( P03DIN )
     ,.P04DIN ( P04DIN ) ,.P05DIN ( P05DIN ) ,.P06DIN ( P06DIN ) ,.P00ENO ( P00ENO )
     ,.P01ENO ( P01ENO ) ,.P02ENO ( P02ENO ) ,.P03ENO ( P03ENO ) ,.P04ENO ( P04ENO )
     ,.P05ENO ( P05ENO ) ,.P06ENO ( P06ENO ) ,.P00PUON ( P00PUON ) ,.P01PUON ( P01PUON )
     ,.P02PUON ( P02PUON ) ,.P03PUON ( P03PUON ) ,.P04PUON ( P04PUON )
     ,.P05PUON ( P05PUON ) ,.P06PUON ( P06PUON ) ,.P00DOUT ( P00DOUT )
     ,.P01DOUT ( P01DOUT ) ,.P02DOUT ( P02DOUT ) ,.P03DOUT ( P03DOUT )
     ,.P04DOUT ( P04DOUT ) ,.P05DOUT ( P05DOUT ) ,.P06DOUT ( P06DOUT )
     ,.P00ENI ( P00ENI ) ,.P01ENI ( P01ENI ) ,.P02ENI ( P02ENI ) ,.P03ENI ( P03ENI )
     ,.P04ENI ( P04ENI ) ,.P05ENI ( P05ENI ) ,.P06ENI ( P06ENI ) ,.PIO00 ( PIO00 )
     ,.PIO01 ( PIO01 ) ,.PIO02 ( PIO02 ) ,.PIO03 ( PIO03 ) ,.PIO04 ( PIO04 )
     ,.PIO05 ( PIO05 ) ,.PIO06 ( PIO06 ) ,.P01SELIN ( P01SELIN ) ,.P03SELIN ( P03SELIN )
     ,.P04SELIN ( P04SELIN ) ,.EXOR ( PORT0EXOR )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_2.0/_macro/_local/kx4_port1v1_mf3_v1.10/_library/100910/kx4_port1v1.hdl
  KX4_PORT1V1 port1 (
    .PCLKRW ( PCLKRW ) ,.PRESETZ ( RESB ) ,.PSEL ( PSELP1 ) ,.PWRITE ( PWRITE )
     ,.PENABLE ( PENABLE ) ,.PADDR4 ( PADDR4 ) ,.PADDR5 ( PADDR5 ) ,.PADDR6 ( PADDR6 )
     ,.PWDATA8 ( MDW8 ) ,.PWDATA9 ( MDW9 ) ,.PWDATA10 ( MDW10 ) ,.PWDATA11 ( MDW11 )
     ,.PWDATA12 ( MDW12 ) ,.PWDATA13 ( MDW13 ) ,.PWDATA14 ( MDW14 ) ,.PWDATA15 ( MDW15 )
     ,.NSRESB ( NSRESB ) ,.SEL64P ( SEL64P ) ,.SEL48P ( SEL48P ) ,.SEL52P ( SEL52P )
     ,.SEL44P ( SEL44P ) ,.SEL36P ( SEL36P ) ,.SEL40P ( SEL40P ) ,.SEL32P ( SEL32P )
     ,.SEL24P ( SEL24P ) ,.SEL08P ( SEL08P ) ,.SEL38P ( SEL38P ) ,.SEL30P ( SEL30P )
     ,.SEL20P ( SEL20P ) ,.SEL64PI ( SEL64PI ) ,.SEL48PI ( SEL48PI ) ,.SEL52PI ( SEL52PI )
     ,.SEL44PI ( SEL44PI ) ,.SEL36PI ( SEL36PI ) ,.SEL40PI ( SEL40PI )
     ,.SEL32PI ( SEL32PI ) ,.SEL24PI ( SEL24PI ) ,.SEL38PI ( SEL38PI )
     ,.SEL30PI ( SEL30PI ) ,.SEL20PI ( SEL20PI ) ,.SCANMODE ( SCANMODE )
     ,.SCANCLK ( SCANCLK ) ,.TESDBT ( TESDBT2 ) ,.OPTOPLRD ( OPTOPLRD )
     ,.PRDATA8 ( PRDP0108 ) ,.PRDATA9 ( PRDP0109 ) ,.PRDATA10 ( PRDP0110 )
     ,.PRDATA11 ( PRDP0111 ) ,.PRDATA12 ( PRDP0112 ) ,.PRDATA13 ( PRDP0113 )
     ,.PRDATA14 ( PRDP0114 ) ,.PRDATA15 ( PRDP0115 ) ,.TESENI0R ( TESENI0R )
     ,.TESENO0R ( TESENO0R ) ,.TDSEL0R ( TDSEL0R ) ,.TDOUT0 ( TDOUT0 )
     ,.TDIN0R ( TDIN0R ) ,.TESENI1R ( TESENI1R ) ,.TESENO1R ( TESENO1R )
     ,.TDSEL1R ( TDSEL1R ) ,.TDOUT1 ( TDOUT1 ) ,.TDIN1R ( TDIN1R ) ,.TESENI2R ( TESENI2R )
     ,.TESENO2R ( TESENO2R ) ,.TDSEL2R ( TDSEL2R ) ,.TDOUT2 ( TDOUT2 )
     ,.TDIN2R ( TDIN2R ) ,.EXINA0 ( P10EXINA ) ,.EXINA1 ( P11EXINA ) ,.EXINA2 ( P12EXINA )
     ,.EXINB0 ( P10EXINB ) ,.EXINA3 ( P13EXINA ) ,.EXINA4 ( P14EXINA )
     ,.EXINB2 ( P12EXINB ) ,.EXINA5 ( P15EXINA ) ,.EXINA6 ( P16EXINA )
     ,.EXINA7 ( P17EXINA ) ,.EXOUTA0 ( P10EXOUTA ) ,.EXOUTA1 ( SOUT010DLY )
     ,.EXOUTA3 ( P13EXOUTA ) ,.EXOUTB1 ( P11EXOUTB ) ,.EXOUTA4 ( SOUT110DLY )
     ,.EXOUTB2 ( P12EXOUTB ) ,.EXOUTC0 ( P10EXOUTC ) ,.EXOUTA5 ( SCKO10 )
     ,.EXOUTB3 ( P13EXOUTB ) ,.EXOUTC1 ( P11EXOUTC ) ,.EXOUTA6 ( P16EXOUTA )
     ,.EXOUTB4 ( P14EXOUTB ) ,.EXOUTC2 ( pull_down72 ) ,.EXOUTA7 ( P17EXOUTA )
     ,.EXOUTB5 ( P15EXOUTB ) ,.EXOUTC3 ( P13EXOUTC ) ,.EXOUTB0 ( P10EXOUTB )
     ,.EXOUTB6 ( TOUT01 ) ,.EXOUTC4 ( P14EXOUTC ) ,.EXOUTB7 ( P17EXOUTB )
     ,.EXOUTC5 ( P15EXOUTC ) ,.EXOUTC6 ( pull_down73 ) ,.EXOUTC7 ( pull_down74 )
     ,.P10DIN ( P10DIN ) ,.P11DIN ( P11DIN ) ,.P12DIN ( P12DIN ) ,.P13DIN ( P13DIN )
     ,.P14DIN ( P14DIN ) ,.P15DIN ( P15DIN ) ,.P16DIN ( P16DIN ) ,.P17DIN ( P17DIN )
     ,.P10ENO ( P10ENO ) ,.P11ENO ( P11ENO ) ,.P12ENO ( P12ENO ) ,.P13ENO ( P13ENO )
     ,.P14ENO ( P14ENO ) ,.P15ENO ( P15ENO ) ,.P16ENO ( P16ENO ) ,.P17ENO ( P17ENO )
     ,.P10PUON ( P10PUON ) ,.P11PUON ( P11PUON ) ,.P12PUON ( P12PUON )
     ,.P13PUON ( P13PUON ) ,.P14PUON ( P14PUON ) ,.P15PUON ( P15PUON )
     ,.P16PUON ( P16PUON ) ,.P17PUON ( P17PUON ) ,.P10DOUT ( P10DOUT )
     ,.P11DOUT ( P11DOUT ) ,.P12DOUT ( P12DOUT ) ,.P13DOUT ( P13DOUT )
     ,.P14DOUT ( P14DOUT ) ,.P15DOUT ( P15DOUT ) ,.P16DOUT ( P16DOUT )
     ,.P17DOUT ( P17DOUT ) ,.P10ENI ( P10ENI ) ,.P11ENI ( P11ENI ) ,.P12ENI ( P12ENI )
     ,.P13ENI ( P13ENI ) ,.P14ENI ( P14ENI ) ,.P15ENI ( P15ENI ) ,.P16ENI ( P16ENI )
     ,.P17ENI ( P17ENI ) ,.PIO10 ( PIO10 ) ,.PIO11 ( PIO11 ) ,.PIO12 ( PIO12 )
     ,.PIO13 ( PIO13 ) ,.PIO14 ( PIO14 ) ,.PIO15 ( PIO15 ) ,.PIO16 ( PIO16 )
     ,.PIO17 ( PIO17 ) ,.P10SELIN ( P10SELIN ) ,.P11SELIN ( P11SELIN )
     ,.P13SELIN ( P13SELIN ) ,.P14SELIN ( P14SELIN ) ,.P15SELIN ( P15SELIN )
     ,.P16SELIN ( P16SELIN ) ,.P17SELIN ( P17SELIN ) ,.TXOCD ( TXOCD )
     ,.TXSAU ( TXSAU ) ,.SLTRXTX ( SLTRXTX ) ,.BBSFDIS1 ( BBSFDIS1 ) ,.EXOR ( PORT1EXOR )
     ,.BBEXAD10 ( BBEXAD10 ) ,.BBEXAD11 ( BBEXAD11 ) ,.BBEXAD12 ( BBEXAD12 )
     ,.BBEXOR10 ( BBEXOR10 ) ,.BBEXOR11 ( BBEXOR11 ) ,.BBEXOR12 ( BBEXOR12 )
     ,.BBMODE ( BBMODE ) ,.BBSWPPT1 ( BBSWPPT1 )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_2.0/_macro/_local/kx4_port2v1_mf3_v1.10/_library/100701/kx4_port2v1.hdl
  KX4_PORT2V1 port2 (
    .PCLKRW ( PCLKRW ) ,.PRESETZ ( RESB ) ,.PSEL ( PSELP2 ) ,.PWRITE ( PWRITE )
     ,.PENABLE ( PENABLE ) ,.PADDR4 ( PADDR4 ) ,.PADDR5 ( PADDR5 ) ,.PADDR6 ( PADDR6 )
     ,.PWDATA0 ( MDW0 ) ,.PWDATA1 ( MDW1 ) ,.PWDATA2 ( MDW2 ) ,.PWDATA3 ( MDW3 )
     ,.PWDATA4 ( MDW4 ) ,.PWDATA5 ( MDW5 ) ,.PWDATA6 ( MDW6 ) ,.PWDATA7 ( MDW7 )
     ,.NSRESB ( NSRESB ) ,.SEL64P ( SEL64P ) ,.SEL48P ( SEL48P ) ,.SEL52P ( SEL52P )
     ,.SEL44P ( SEL44P ) ,.SEL36P ( SEL36P ) ,.SEL40P ( SEL40P ) ,.SEL32P ( SEL32P )
     ,.SEL24P ( SEL24P ) ,.SEL08P ( SEL08P ) ,.SEL38P ( SEL38P ) ,.SEL30P ( SEL30P )
     ,.SEL20P ( SEL20P ) ,.SEL64PI ( SEL64PI ) ,.SEL48PI ( SEL48PI ) ,.SEL52PI ( SEL52PI )
     ,.SEL44PI ( SEL44PI ) ,.SEL36PI ( SEL36PI ) ,.SEL40PI ( SEL40PI )
     ,.SEL32PI ( SEL32PI ) ,.SEL24PI ( SEL24PI ) ,.SEL38PI ( SEL38PI )
     ,.SEL30PI ( SEL30PI ) ,.SEL20PI ( SEL20PI ) ,.SCANMODE ( SCANMODE )
     ,.SCANCLK ( SCANCLK ) ,.TESDBT ( TESDBT2 ) ,.OPTOPLRD ( OPTOPLRD )
     ,.TESENO0T ( TESENO0T ) ,.TESENO1T ( TESENO1T ) ,.TESENO2T ( TESENO2T )
     ,.TESENI0T ( TESENI0T ) ,.TESENI1T ( TESENI1T ) ,.TESENI2T ( TESENI2T )
     ,.TDSEL0T ( TDSEL0T ) ,.TDSEL1T ( TDSEL1T ) ,.TDSEL2T ( TDSEL2T )
     ,.TDOUT0 ( TDOUT0 ) ,.TDOUT1 ( TDOUT1 ) ,.TDOUT2 ( TDOUT2 ) ,.TDIN0T ( TDIN0T )
     ,.TDIN1T ( TDIN1T ) ,.TDIN2T ( TDIN2T ) ,.PRDATA0 ( PRDP0200 ) ,.PRDATA1 ( PRDP0201 )
     ,.PRDATA2 ( PRDP0202 ) ,.PRDATA3 ( PRDP0203 ) ,.PRDATA4 ( PRDP0204 )
     ,.PRDATA5 ( PRDP0205 ) ,.PRDATA6 ( PRDP0206 ) ,.PRDATA7 ( PRDP0207 )
     ,.DGEN00 ( DGEN00 ) ,.DGEN01 ( DGEN01 ) ,.DGEN02 ( DGEN02 ) ,.DGEN03 ( DGEN03 )
     ,.DGEN04 ( DGEN04 ) ,.DGEN05 ( DGEN05 ) ,.DGEN06 ( DGEN06 ) ,.DGEN07 ( DGEN07 )
     ,.P20DIN ( P20DIN ) ,.P21DIN ( P21DIN ) ,.P22DIN ( P22DIN ) ,.P23DIN ( P23DIN )
     ,.P24DIN ( P24DIN ) ,.P25DIN ( P25DIN ) ,.P26DIN ( P26DIN ) ,.P27DIN ( P27DIN )
     ,.P20ENO ( P20ENO ) ,.P21ENO ( P21ENO ) ,.P22ENO ( P22ENO ) ,.P23ENO ( P23ENO )
     ,.P24ENO ( P24ENO ) ,.P25ENO ( P25ENO ) ,.P26ENO ( P26ENO ) ,.P27ENO ( P27ENO )
     ,.P20DOUT ( P20DOUT ) ,.P21DOUT ( P21DOUT ) ,.P22DOUT ( P22DOUT )
     ,.P23DOUT ( P23DOUT ) ,.P24DOUT ( P24DOUT ) ,.P25DOUT ( P25DOUT )
     ,.P26DOUT ( P26DOUT ) ,.P27DOUT ( P27DOUT ) ,.P20ENI ( P20ENI ) ,.P21ENI ( P21ENI )
     ,.P22ENI ( P22ENI ) ,.P23ENI ( P23ENI ) ,.P24ENI ( P24ENI ) ,.P25ENI ( P25ENI )
     ,.P26ENI ( P26ENI ) ,.P27ENI ( P27ENI ) ,.PIO20 ( PIO20 ) ,.PIO21 ( PIO21 )
     ,.PIO22 ( PIO22 ) ,.PIO23 ( PIO23 ) ,.PIO24 ( PIO24 ) ,.PIO25 ( PIO25 )
     ,.PIO26 ( PIO26 ) ,.PIO27 ( PIO27 ) ,.EXOR ( PORT2EXOR )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_2.0/_macro/_local/kx4_port3v1_mf3_v1.10/_library/100701/kx4_port3v1.hdl
  KX4_PORT3V1 port3 (
    .PCLKRW ( PCLKRW ) ,.PRESETZ ( RESB ) ,.PSEL ( PSELP3 ) ,.PWRITE ( PWRITE )
     ,.PENABLE ( PENABLE ) ,.PADDR4 ( PADDR4 ) ,.PADDR5 ( PADDR5 ) ,.PADDR6 ( PADDR6 )
     ,.PWDATA8 ( MDW8 ) ,.PWDATA9 ( MDW9 ) ,.NSRESB ( NSRESB ) ,.SEL64P ( SEL64P )
     ,.SEL48P ( SEL48P ) ,.SEL52P ( SEL52P ) ,.SEL44P ( SEL44P ) ,.SEL36P ( SEL36P )
     ,.SEL40P ( SEL40P ) ,.SEL32P ( SEL32P ) ,.SEL24P ( SEL24P ) ,.SEL08P ( SEL08P )
     ,.SEL38P ( SEL38P ) ,.SEL30P ( SEL30P ) ,.SEL20P ( SEL20P ) ,.SEL64PI ( SEL64PI )
     ,.SEL48PI ( SEL48PI ) ,.SEL52PI ( SEL52PI ) ,.SEL44PI ( SEL44PI )
     ,.SEL36PI ( SEL36PI ) ,.SEL40PI ( SEL40PI ) ,.SEL32PI ( SEL32PI )
     ,.SEL24PI ( SEL24PI ) ,.SEL38PI ( SEL38PI ) ,.SEL30PI ( SEL30PI )
     ,.SEL20PI ( SEL20PI ) ,.SCANMODE ( SCANMODE ) ,.SCANCLK ( SCANCLK )
     ,.TESDBT ( TESDBT2 ) ,.OPTOPLRD ( OPTOPLRD ) ,.PRDATA8 ( PRDP0308 )
     ,.PRDATA9 ( PRDP0309 ) ,.PRDATA10 ( PRDP0310 ) ,.PRDATA11 ( PRDP0311 )
     ,.PRDATA12 ( PRDP0312 ) ,.PRDATA13 ( PRDP0313 ) ,.PRDATA14 ( PRDP0314 )
     ,.PRDATA15 ( PRDP0315 ) ,.EXINA0 ( P30EXINA ) ,.EXINA1 ( P31EXINA )
     ,.EXOUTA0 ( SCKO03 ) ,.EXOUTA1 ( pull_up63 ) ,.EXOUTB0 ( CLK1HZ )
     ,.EXOUTB1 ( P31EXOUTB ) ,.EXOUTC0 ( pull_down75 ) ,.EXOUTC1 ( P31EXOUTC )
     ,.P30DIN ( P30DIN ) ,.P31DIN ( P31DIN ) ,.P30ENO ( P30ENO ) ,.P31ENO ( P31ENO )
     ,.P30PUON ( P30PUON ) ,.P31PUON ( P31PUON ) ,.P30DOUT ( P30DOUT )
     ,.P31DOUT ( P31DOUT ) ,.P30ENI ( P30ENI ) ,.P31ENI ( P31ENI ) ,.PIO30 ( PIO30 )
     ,.PIO31 ( PIO31 ) ,.EXOR ( PORT3EXOR )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_2.0/_macro/_local/kx4_port4v1_mf3_v1.10/_library/100701/kx4_port4v1.hdl
  KX4_PORT4V1 port4 (
    .PCLKRW ( PCLKRW ) ,.PRESETZ ( RESB ) ,.PSEL ( PSELP4 ) ,.PWRITE ( PWRITE )
     ,.PENABLE ( PENABLE ) ,.PADDR4 ( PADDR4 ) ,.PADDR5 ( PADDR5 ) ,.PADDR6 ( PADDR6 )
     ,.PWDATA0 ( MDW0 ) ,.PWDATA1 ( MDW1 ) ,.PWDATA2 ( MDW2 ) ,.PWDATA3 ( MDW3 )
     ,.NSRESB ( NSRESB ) ,.SEL64P ( SEL64P ) ,.SEL48P ( SEL48P ) ,.SEL52P ( SEL52P )
     ,.SEL44P ( SEL44P ) ,.SEL36P ( SEL36P ) ,.SEL40P ( SEL40P ) ,.SEL32P ( SEL32P )
     ,.SEL24P ( SEL24P ) ,.SEL08P ( SEL08P ) ,.SEL38P ( SEL38P ) ,.SEL30P ( SEL30P )
     ,.SEL20P ( SEL20P ) ,.SEL64PI ( SEL64PI ) ,.SEL48PI ( SEL48PI ) ,.SEL52PI ( SEL52PI )
     ,.SEL44PI ( SEL44PI ) ,.SEL36PI ( SEL36PI ) ,.SEL40PI ( SEL40PI )
     ,.SEL32PI ( SEL32PI ) ,.SEL24PI ( SEL24PI ) ,.SEL38PI ( SEL38PI )
     ,.SEL30PI ( SEL30PI ) ,.SEL20PI ( SEL20PI ) ,.SCANMODE ( SCANMODE )
     ,.SCANCLK ( SCANCLK ) ,.TESDBT ( TESDBT2 ) ,.OPTOPLRD ( OPTOPLRD )
     ,.TSELOREG ( TSELOREG ) ,.TSELIRES ( TSELIRES ) ,.TTEMP ( TTEMP )
     ,.TESENO3 ( TESENO3 ) ,.TESENI3 ( TESENI3 ) ,.TDSEL3 ( TDSEL3 ) ,.TDOUT3 ( TDOUT3 )
     ,.TDIN3 ( TDIN3 ) ,.PRDATA0 ( PRDP0400 ) ,.PRDATA1 ( PRDP0401 ) ,.PRDATA2 ( PRDP0402 )
     ,.PRDATA3 ( PRDP0403 ) ,.PRDATA4 ( PRDP0404 ) ,.PRDATA5 ( PRDP0405 )
     ,.PRDATA6 ( PRDP0406 ) ,.PRDATA7 ( PRDP0407 ) ,.RXOCD ( RXOCD ) ,.EXINA1 ( P41EXINA )
     ,.EXINA2 ( P42EXINA ) ,.EXINA3 ( P43EXINA ) ,.TXOCD ( TXOCD ) ,.EXOUTA1 ( pull_up64 )
     ,.EXOUTA2 ( pull_up65 ) ,.EXOUTA3 ( pull_up66 ) ,.EXOUTB1 ( P41EXOUTB )
     ,.EXOUTB2 ( P42EXOUTB ) ,.EXOUTB3 ( pull_down78 ) ,.EXOUTC1 ( pull_down76 )
     ,.EXOUTC2 ( pull_down77 ) ,.EXOUTC3 ( pull_down79 ) ,.OCDMOD ( OCDMOD )
     ,.SPRGMOD ( SPRGMOD ) ,.GOFIRM ( GOFIRM ) ,.SLTRXTX ( SLTRXTX ) ,.P40DIN ( P40DIN )
     ,.P41DIN ( P41DIN ) ,.P42DIN ( P42DIN ) ,.P43DIN ( P43DIN ) ,.P40ENO ( P40ENO )
     ,.P41ENO ( P41ENO ) ,.P42ENO ( P42ENO ) ,.P43ENO ( P43ENO ) ,.P40PUON ( P40PUON )
     ,.P41PUON ( P41PUON ) ,.P42PUON ( P42PUON ) ,.P43PUON ( P43PUON )
     ,.P40DOUT ( P40DOUT ) ,.P41DOUT ( P41DOUT ) ,.P42DOUT ( P42DOUT )
     ,.P43DOUT ( P43DOUT ) ,.P40ENI ( P40ENI ) ,.P41ENI ( P41ENI ) ,.P42ENI ( P42ENI )
     ,.P43ENI ( P43ENI ) ,.PIO40 ( PIO40 ) ,.PIO41 ( PIO41 ) ,.PIO42 ( PIO42 )
     ,.PIO43 ( PIO43 ) ,.EXOR ( PORT4EXOR )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_2.0/_macro/_local/kx4_port5v1_mf3_v1.10/_library/100701/kx4_port5v1.hdl
  KX4_PORT5V1 port5 (
    .PCLKRW ( PCLKRW ) ,.PRESETZ ( RESB ) ,.PSEL ( PSELP5 ) ,.PWRITE ( PWRITE )
     ,.PENABLE ( PENABLE ) ,.PADDR4 ( PADDR4 ) ,.PADDR5 ( PADDR5 ) ,.PADDR6 ( PADDR6 )
     ,.PWDATA8 ( MDW8 ) ,.PWDATA9 ( MDW9 ) ,.PWDATA10 ( MDW10 ) ,.PWDATA11 ( MDW11 )
     ,.PWDATA12 ( MDW12 ) ,.PWDATA13 ( MDW13 ) ,.NSRESB ( NSRESB ) ,.SEL64P ( SEL64P )
     ,.SEL48P ( SEL48P ) ,.SEL52P ( SEL52P ) ,.SEL44P ( SEL44P ) ,.SEL36P ( SEL36P )
     ,.SEL40P ( SEL40P ) ,.SEL32P ( SEL32P ) ,.SEL24P ( SEL24P ) ,.SEL08P ( SEL08P )
     ,.SEL38P ( SEL38P ) ,.SEL30P ( SEL30P ) ,.SEL20P ( SEL20P ) ,.SEL64PI ( SEL64PI )
     ,.SEL48PI ( SEL48PI ) ,.SEL52PI ( SEL52PI ) ,.SEL44PI ( SEL44PI )
     ,.SEL36PI ( SEL36PI ) ,.SEL40PI ( SEL40PI ) ,.SEL32PI ( SEL32PI )
     ,.SEL24PI ( SEL24PI ) ,.SEL38PI ( SEL38PI ) ,.SEL30PI ( SEL30PI )
     ,.SEL20PI ( SEL20PI ) ,.SCANMODE ( SCANMODE ) ,.SCANCLK ( SCANCLK )
     ,.TESDBT ( TESDBT2 ) ,.OPTOPLRD ( OPTOPLRD ) ,.PRDATA8 ( PRDP0508 )
     ,.PRDATA9 ( PRDP0509 ) ,.PRDATA10 ( PRDP0510 ) ,.PRDATA11 ( PRDP0511 )
     ,.PRDATA12 ( PRDP0512 ) ,.PRDATA13 ( PRDP0513 ) ,.PRDATA14 ( PRDP0514 )
     ,.PRDATA15 ( PRDP0515 ) ,.EXINA0 ( P50EXINA ) ,.EXINA1 ( P51EXINA )
     ,.EXINA2 ( P52EXINA ) ,.EXINA3 ( P53EXINA ) ,.EXINA4 ( P54EXINA )
     ,.EXINA5 ( P55EXINA ) ,.EXOUTA0 ( SOUT013DLY ) ,.EXOUTA1 ( P51EXOUTA )
     ,.EXOUTA2 ( pull_up67 ) ,.EXOUTB0 ( pull_down80 ) ,.EXOUTA3 ( pull_up68 )
     ,.EXOUTB1 ( pull_down82 ) ,.EXOUTA4 ( pull_up69 ) ,.EXOUTB2 ( pull_down84 )
     ,.EXOUTC0 ( pull_down81 ) ,.EXOUTA5 ( P55EXOUTA ) ,.EXOUTB3 ( pull_down86 )
     ,.EXOUTC1 ( pull_down83 ) ,.EXOUTB4 ( pull_down88 ) ,.EXOUTC2 ( pull_down85 )
     ,.EXOUTB5 ( P55EXOUTB ) ,.EXOUTC3 ( pull_down87 ) ,.EXOUTC4 ( pull_down89 )
     ,.EXOUTC5 ( pull_down90 ) ,.P50DIN ( P50DIN ) ,.P51DIN ( P51DIN )
     ,.P52DIN ( P52DIN ) ,.P53DIN ( P53DIN ) ,.P54DIN ( P54DIN ) ,.P55DIN ( P55DIN )
     ,.P50ENO ( P50ENO ) ,.P51ENO ( P51ENO ) ,.P52ENO ( P52ENO ) ,.P53ENO ( P53ENO )
     ,.P54ENO ( P54ENO ) ,.P55ENO ( P55ENO ) ,.P50PUON ( P50PUON ) ,.P51PUON ( P51PUON )
     ,.P52PUON ( P52PUON ) ,.P53PUON ( P53PUON ) ,.P54PUON ( P54PUON )
     ,.P55PUON ( P55PUON ) ,.P50DOUT ( P50DOUT ) ,.P51DOUT ( P51DOUT )
     ,.P52DOUT ( P52DOUT ) ,.P53DOUT ( P53DOUT ) ,.P54DOUT ( P54DOUT )
     ,.P55DOUT ( P55DOUT ) ,.P50ENI ( P50ENI ) ,.P51ENI ( P51ENI ) ,.P52ENI ( P52ENI )
     ,.P53ENI ( P53ENI ) ,.P54ENI ( P54ENI ) ,.P55ENI ( P55ENI ) ,.PIO50 ( PIO50 )
     ,.PIO51 ( PIO51 ) ,.PIO52 ( PIO52 ) ,.PIO53 ( PIO53 ) ,.PIO54 ( PIO54 )
     ,.PIO55 ( PIO55 ) ,.P55SELIN ( P55SELIN ) ,.EXOR ( PORT5EXOR )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_2.0/_macro/_local/kx4_port6v1_mf3_v1.10/_library/100701/kx4_port6v1.hdl
  KX4_PORT6V1 port6 (
    .PCLKRW ( PCLKRW ) ,.PRESETZ ( RESB ) ,.PSEL ( PSELP6 ) ,.PWRITE ( PWRITE )
     ,.PENABLE ( PENABLE ) ,.PADDR4 ( PADDR4 ) ,.PADDR5 ( PADDR5 ) ,.PADDR6 ( PADDR6 )
     ,.PWDATA0 ( MDW0 ) ,.PWDATA1 ( MDW1 ) ,.PWDATA2 ( MDW2 ) ,.PWDATA3 ( MDW3 )
     ,.NSRESB ( NSRESB ) ,.SEL64P ( SEL64P ) ,.SEL48P ( SEL48P ) ,.SEL52P ( SEL52P )
     ,.SEL44P ( SEL44P ) ,.SEL36P ( SEL36P ) ,.SEL40P ( SEL40P ) ,.SEL32P ( SEL32P )
     ,.SEL24P ( SEL24P ) ,.SEL08P ( SEL08P ) ,.SEL38P ( SEL38P ) ,.SEL30P ( SEL30P )
     ,.SEL20P ( SEL20P ) ,.SEL64PI ( SEL64PI ) ,.SEL48PI ( SEL48PI ) ,.SEL52PI ( SEL52PI )
     ,.SEL44PI ( SEL44PI ) ,.SEL36PI ( SEL36PI ) ,.SEL40PI ( SEL40PI )
     ,.SEL32PI ( SEL32PI ) ,.SEL24PI ( SEL24PI ) ,.SEL38PI ( SEL38PI )
     ,.SEL30PI ( SEL30PI ) ,.SEL20PI ( SEL20PI ) ,.SCANMODE ( SCANMODE )
     ,.SCANCLK ( SCANCLK ) ,.TESDBT ( TESDBT2 ) ,.OPTOPLRD ( OPTOPLRD )
     ,.PRDATA0 ( PRDP0600 ) ,.PRDATA1 ( PRDP0601 ) ,.PRDATA2 ( PRDP0602 )
     ,.PRDATA3 ( PRDP0603 ) ,.PRDATA4 ( PRDP0604 ) ,.PRDATA5 ( PRDP0605 )
     ,.PRDATA6 ( PRDP0606 ) ,.PRDATA7 ( PRDP0607 ) ,.EXINA0 ( P60EXINA )
     ,.EXINA1 ( P61EXINA ) ,.EXINA2 ( P62EXINA ) ,.EXINA3 ( P63EXINA )
     ,.EXOUTA0 ( pull_up70 ) ,.EXOUTA1 ( pull_up71 ) ,.EXOUTA2 ( pull_up72 )
     ,.EXOUTB0 ( P60EXOUTB ) ,.EXOUTA3 ( pull_up73 ) ,.EXOUTB1 ( P61EXOUTB )
     ,.EXOUTB2 ( pull_down93 ) ,.EXOUTC0 ( pull_down91 ) ,.EXOUTB3 ( pull_down95 )
     ,.EXOUTC1 ( pull_down92 ) ,.EXOUTC2 ( pull_down94 ) ,.EXOUTC3 ( pull_down96 )
     ,.P60DIN ( P60DIN ) ,.P61DIN ( P61DIN ) ,.P62DIN ( P62DIN ) ,.P63DIN ( P63DIN )
     ,.P60ENO ( P60ENO ) ,.P61ENO ( P61ENO ) ,.P62ENO ( P62ENO ) ,.P63ENO ( P63ENO )
     ,.P60DOUT ( P60DOUT ) ,.P61DOUT ( P61DOUT ) ,.P62DOUT ( P62DOUT )
     ,.P63DOUT ( P63DOUT ) ,.P60ENI ( P60ENI ) ,.P61ENI ( P61ENI ) ,.P62ENI ( P62ENI )
     ,.P63ENI ( P63ENI ) ,.PIO60 ( PIO60 ) ,.PIO61 ( PIO61 ) ,.PIO62 ( PIO62 )
     ,.PIO63 ( PIO63 ) ,.EXOR ( PORT6EXOR )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_2.0/_macro/_local/kx4_port7v1_mf3_v1.10/_library/100701/kx4_port7v1.hdl
  KX4_PORT7V1 port7 (
    .PCLKRW ( PCLKRW ) ,.PRESETZ ( RESB ) ,.PSEL ( PSELP7 ) ,.PWRITE ( PWRITE )
     ,.PENABLE ( PENABLE ) ,.PADDR4 ( PADDR4 ) ,.PADDR5 ( PADDR5 ) ,.PADDR6 ( PADDR6 )
     ,.PWDATA8 ( MDW8 ) ,.PWDATA9 ( MDW9 ) ,.PWDATA10 ( MDW10 ) ,.PWDATA11 ( MDW11 )
     ,.PWDATA12 ( MDW12 ) ,.PWDATA13 ( MDW13 ) ,.PWDATA14 ( MDW14 ) ,.PWDATA15 ( MDW15 )
     ,.NSRESB ( NSRESB ) ,.PSELKR ( PSELKR ) ,.INTKR ( INTKR ) ,.SEL64P ( SEL64P )
     ,.SEL48P ( SEL48P ) ,.SEL52P ( SEL52P ) ,.SEL44P ( SEL44P ) ,.SEL36P ( SEL36P )
     ,.SEL40P ( SEL40P ) ,.SEL32P ( SEL32P ) ,.SEL24P ( SEL24P ) ,.SEL08P ( SEL08P )
     ,.SEL38P ( SEL38P ) ,.SEL30P ( SEL30P ) ,.SEL20P ( SEL20P ) ,.SEL64PI ( SEL64PI )
     ,.SEL48PI ( SEL48PI ) ,.SEL52PI ( SEL52PI ) ,.SEL44PI ( SEL44PI )
     ,.SEL36PI ( SEL36PI ) ,.SEL40PI ( SEL40PI ) ,.SEL32PI ( SEL32PI )
     ,.SEL24PI ( SEL24PI ) ,.SEL38PI ( SEL38PI ) ,.SEL30PI ( SEL30PI )
     ,.SEL20PI ( SEL20PI ) ,.SCANMODE ( SCANMODE ) ,.SCANCLK ( SCANCLK )
     ,.TESDBT ( TESDBT2 ) ,.OPTOPLRD ( OPTOPLRD ) ,.PRDATA8 ( PRDP0708 )
     ,.PRDATA9 ( PRDP0709 ) ,.PRDATA10 ( PRDP0710 ) ,.PRDATA11 ( PRDP0711 )
     ,.PRDATA12 ( PRDP0712 ) ,.PRDATA13 ( PRDP0713 ) ,.PRDATA14 ( PRDP0714 )
     ,.PRDATA15 ( PRDP0715 ) ,.TESENI0B ( TESENI0B ) ,.TESENO0B ( TESENO0B )
     ,.TDSEL0B ( TDSEL0B ) ,.TDOUT0 ( TDOUT0 ) ,.TDIN0B ( TDIN0B ) ,.TESENI1B ( TESENI1B )
     ,.TESENO1B ( TESENO1B ) ,.TDSEL1B ( TDSEL1B ) ,.TDOUT1 ( TDOUT1 )
     ,.TDIN1B ( TDIN1B ) ,.TESENI2B ( TESENI2B ) ,.TESENO2B ( TESENO2B )
     ,.TDSEL2B ( TDSEL2B ) ,.TDOUT2 ( TDOUT2 ) ,.TDIN2B ( TDIN2B ) ,.EXINA0 ( P70EXINA )
     ,.EXINA1 ( P71EXINA ) ,.EXINA2 ( P72EXINA ) ,.EXINA3 ( P73EXINA )
     ,.EXINA4 ( P74EXINA ) ,.EXINA5 ( P75EXINA ) ,.EXINA6 ( P76EXINA )
     ,.EXINA7 ( P77EXINA ) ,.EXOUTA0 ( SCKO11 ) ,.EXOUTA1 ( SOUT111DLY )
     ,.EXOUTA2 ( SOUT101 ) ,.EXOUTB0 ( pull_down97 ) ,.EXOUTA3 ( SOUT001 )
     ,.EXOUTB1 ( pull_down99 ) ,.EXOUTA4 ( SOUT011DLY ) ,.EXOUTB2 ( pull_down101 )
     ,.EXOUTC0 ( pull_down98 ) ,.EXOUTA5 ( SCKO01 ) ,.EXOUTB3 ( pull_down103 )
     ,.EXOUTC1 ( pull_down100 ) ,.EXOUTA6 ( pull_up74 ) ,.EXOUTB4 ( pull_down105 )
     ,.EXOUTC2 ( pull_down102 ) ,.EXOUTA7 ( P77EXOUTA ) ,.EXOUTB5 ( pull_down107 )
     ,.EXOUTC3 ( pull_down104 ) ,.EXOUTB6 ( pull_down109 ) ,.EXOUTC4 ( pull_down106 )
     ,.EXOUTB7 ( pull_down111 ) ,.EXOUTC5 ( pull_down108 ) ,.EXOUTC6 ( pull_down110 )
     ,.EXOUTC7 ( pull_down112 ) ,.P70DIN ( P70DIN ) ,.P71DIN ( P71DIN )
     ,.P72DIN ( P72DIN ) ,.P73DIN ( P73DIN ) ,.P74DIN ( P74DIN ) ,.P75DIN ( P75DIN )
     ,.P76DIN ( P76DIN ) ,.P77DIN ( P77DIN ) ,.P70ENO ( P70ENO ) ,.P71ENO ( P71ENO )
     ,.P72ENO ( P72ENO ) ,.P73ENO ( P73ENO ) ,.P74ENO ( P74ENO ) ,.P75ENO ( P75ENO )
     ,.P76ENO ( P76ENO ) ,.P77ENO ( P77ENO ) ,.P70PUON ( P70PUON ) ,.P71PUON ( P71PUON )
     ,.P72PUON ( P72PUON ) ,.P73PUON ( P73PUON ) ,.P74PUON ( P74PUON )
     ,.P75PUON ( P75PUON ) ,.P76PUON ( P76PUON ) ,.P77PUON ( P77PUON )
     ,.P70DOUT ( P70DOUT ) ,.P71DOUT ( P71DOUT ) ,.P72DOUT ( P72DOUT )
     ,.P73DOUT ( P73DOUT ) ,.P74DOUT ( P74DOUT ) ,.P75DOUT ( P75DOUT )
     ,.P76DOUT ( P76DOUT ) ,.P77DOUT ( P77DOUT ) ,.P70ENI ( P70ENI ) ,.P71ENI ( P71ENI )
     ,.P72ENI ( P72ENI ) ,.P73ENI ( P73ENI ) ,.P74ENI ( P74ENI ) ,.P75ENI ( P75ENI )
     ,.P76ENI ( P76ENI ) ,.P77ENI ( P77ENI ) ,.PIO70 ( PIO70 ) ,.PIO71 ( PIO71 )
     ,.PIO72 ( PIO72 ) ,.PIO73 ( PIO73 ) ,.PIO74 ( PIO74 ) ,.PIO75 ( PIO75 )
     ,.PIO76 ( PIO76 ) ,.PIO77 ( PIO77 ) ,.CLK60MHZ ( CLK60MHZ ) ,.EXOR ( PORT7EXOR )
    
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_2.0/_macro/_local/kx4_port12v1_mf3_v1.10/_library/100701/kx4_port12v1.hdl
  KX4_PORT12V1 port12 (
    .PCLKRW ( PCLKRW ) ,.PRESETZ ( RESB ) ,.PSEL ( PSELP12 ) ,.PWRITE ( PWRITE )
     ,.PENABLE ( PENABLE ) ,.PADDR4 ( PADDR4 ) ,.PADDR5 ( PADDR5 ) ,.PADDR6 ( PADDR6 )
     ,.PWDATA0 ( MDW0 ) ,.NSRESB ( NSRESB ) ,.SEL64P ( SEL64P ) ,.SEL48P ( SEL48P )
     ,.SEL52P ( SEL52P ) ,.SEL44P ( SEL44P ) ,.SEL36P ( SEL36P ) ,.SEL40P ( SEL40P )
     ,.SEL32P ( SEL32P ) ,.SEL24P ( SEL24P ) ,.SEL08P ( SEL08P ) ,.SEL38P ( SEL38P )
     ,.SEL30P ( SEL30P ) ,.SEL20P ( SEL20P ) ,.SEL64PI ( SEL64PI ) ,.SEL48PI ( SEL48PI )
     ,.SEL52PI ( SEL52PI ) ,.SEL44PI ( SEL44PI ) ,.SEL36PI ( SEL36PI )
     ,.SEL40PI ( SEL40PI ) ,.SEL32PI ( SEL32PI ) ,.SEL24PI ( SEL24PI )
     ,.SEL38PI ( SEL38PI ) ,.SEL30PI ( SEL30PI ) ,.SEL20PI ( SEL20PI )
     ,.SCANMODE ( SCANMODE ) ,.SCANCLK ( SCANCLK ) ,.TESDBT ( TESDBT2 )
     ,.OPTOPLRD ( OPTOPLRD ) ,.TESENI4 ( TESENI4 ) ,.TDIN4 ( TDIN4 ) ,.PRDATA0 ( PRDP1200 )
     ,.PRDATA1 ( PRDP1201 ) ,.PRDATA2 ( PRDP1202 ) ,.PRDATA3 ( PRDP1203 )
     ,.PRDATA4 ( PRDP1204 ) ,.PRDATA5 ( PRDP1205 ) ,.PRDATA6 ( PRDP1206 )
     ,.PRDATA7 ( PRDP1207 ) ,.EXINA0 ( P120EXINA ) ,.EXINA2 ( P122EXINA )
     ,.EXOUTA0 ( pull_up75 ) ,.EXOUTB0 ( pull_down113 ) ,.EXOUTC0 ( pull_down114 )
     ,.P120DIN ( P120DIN ) ,.P121DIN ( X1DIN ) ,.P122DIN ( X2DIN ) ,.P123DIN ( XT1DIN )
     ,.P124DIN ( XT2DIN ) ,.P120ENO ( P120ENO ) ,.P120PUON ( P120PUON )
     ,.P120DOUT ( P120DOUT ) ,.P120ENI ( P120ENI ) ,.P121ENI ( X1ENI )
     ,.P122ENI ( X2ENI ) ,.P123ENI ( XT1ENI ) ,.P124ENI ( XT2ENI ) ,.PIO120 ( PIO120 )
     ,.PIO121 ( PIO121 ) ,.PIO122 ( PIO122 ) ,.PIO123 ( PIO123 ) ,.PIO124 ( PIO124 )
     ,.EXOR ( PORT12EXOR )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_2.0/_macro/_local/kx4_port13v1_mf3_v1.10/_library/100904/kx4_port13v1.hdl
  KX4_PORT13V1 port13 (
    .PCLKRW ( PCLKRW ) ,.PRESETZ ( RESB ) ,.PSEL ( PSELP13 ) ,.PWRITE ( PWRITE )
     ,.PENABLE ( PENABLE ) ,.PADDR4 ( PADDR4 ) ,.PADDR5 ( PADDR5 ) ,.PADDR6 ( PADDR6 )
     ,.PWDATA8 ( MDW8 ) ,.NSRESB ( NSRESB ) ,.SEL64P ( SEL64P ) ,.SEL48P ( SEL48P )
     ,.SEL52P ( SEL52P ) ,.SEL44P ( SEL44P ) ,.SEL36P ( SEL36P ) ,.SEL40P ( SEL40P )
     ,.SEL32P ( SEL32P ) ,.SEL24P ( SEL24P ) ,.SEL08P ( SEL08P ) ,.SEL38P ( SEL38P )
     ,.SEL30P ( SEL30P ) ,.SEL20P ( SEL20P ) ,.SEL64PI ( SEL64PI ) ,.SEL48PI ( SEL48PI )
     ,.SEL52PI ( SEL52PI ) ,.SEL44PI ( SEL44PI ) ,.SEL36PI ( SEL36PI )
     ,.SEL40PI ( SEL40PI ) ,.SEL32PI ( SEL32PI ) ,.SEL24PI ( SEL24PI )
     ,.SEL38PI ( SEL38PI ) ,.SEL30PI ( SEL30PI ) ,.SEL20PI ( SEL20PI )
     ,.SCANMODE ( SCANMODE ) ,.TESDBT ( TESDBT2 ) ,.TDIN5 ( TDIN5 ) ,.PRDATA8 ( PRDP1308 )
     ,.PRDATA9 ( PRDP1309 ) ,.PRDATA10 ( PRDP1310 ) ,.PRDATA11 ( PRDP1311 )
     ,.PRDATA12 ( PRDP1312 ) ,.PRDATA13 ( PRDP1313 ) ,.PRDATA14 ( PRDP1314 )
     ,.PRDATA15 ( PRDP1315 ) ,.MODIDIS ( MODIDIS ) ,.EXINA7 ( P137EXINA )
     ,.P137DIN ( P137DIN ) ,.P130ENO ( P130ENO ) ,.P130DOUT ( P130DOUT )
     ,.P137ENI ( P137ENI ) ,.PIO130 ( PIO130 ) ,.PIO137 ( PIO137 )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_2.0/_macro/_local/kx4_port14v1_mf3_v1.10/_library/100701/kx4_port14v1.hdl
  KX4_PORT14V1 port14 (
    .PCLKRW ( PCLKRW ) ,.PRESETZ ( RESB ) ,.PSEL ( PSELP14 ) ,.PWRITE ( PWRITE )
     ,.PENABLE ( PENABLE ) ,.PADDR4 ( PADDR4 ) ,.PADDR5 ( PADDR5 ) ,.PADDR6 ( PADDR6 )
     ,.PWDATA0 ( MDW0 ) ,.PWDATA1 ( MDW1 ) ,.PWDATA6 ( MDW6 ) ,.PWDATA7 ( MDW7 )
     ,.NSRESB ( NSRESB ) ,.SEL64P ( SEL64P ) ,.SEL48P ( SEL48P ) ,.SEL52P ( SEL52P )
     ,.SEL44P ( SEL44P ) ,.SEL36P ( SEL36P ) ,.SEL40P ( SEL40P ) ,.SEL32P ( SEL32P )
     ,.SEL24P ( SEL24P ) ,.SEL08P ( SEL08P ) ,.SEL38P ( SEL38P ) ,.SEL30P ( SEL30P )
     ,.SEL20P ( SEL20P ) ,.SEL64PI ( SEL64PI ) ,.SEL48PI ( SEL48PI ) ,.SEL52PI ( SEL52PI )
     ,.SEL44PI ( SEL44PI ) ,.SEL36PI ( SEL36PI ) ,.SEL40PI ( SEL40PI )
     ,.SEL32PI ( SEL32PI ) ,.SEL24PI ( SEL24PI ) ,.SEL38PI ( SEL38PI )
     ,.SEL30PI ( SEL30PI ) ,.SEL20PI ( SEL20PI ) ,.SCANMODE ( SCANMODE )
     ,.SCANCLK ( SCANCLK ) ,.TESDBT ( TESDBT2 ) ,.OPTOPLRD ( OPTOPLRD )
     ,.PRDATA0 ( PRDP1400 ) ,.PRDATA1 ( PRDP1401 ) ,.PRDATA2 ( PRDP1402 )
     ,.PRDATA3 ( PRDP1403 ) ,.PRDATA4 ( PRDP1404 ) ,.PRDATA5 ( PRDP1405 )
     ,.PRDATA6 ( PRDP1406 ) ,.PRDATA7 ( PRDP1407 ) ,.EXINA0 ( P140EXINA )
     ,.EXINA1 ( P141EXINA ) ,.EXINA6 ( P146EXINA ) ,.EXINA7 ( P147EXINA )
     ,.EXOUTA0 ( pull_up76 ) ,.EXOUTA1 ( pull_up77 ) ,.EXOUTA6 ( pull_up78 )
     ,.EXOUTA7 ( pull_up79 ) ,.EXOUTB0 ( P140EXOUTB ) ,.EXOUTB1 ( P141EXOUTB )
     ,.EXOUTB6 ( pull_down117 ) ,.EXOUTB7 ( pull_down119 ) ,.EXOUTC0 ( pull_down115 )
     ,.EXOUTC1 ( pull_down116 ) ,.EXOUTC6 ( pull_down118 ) ,.EXOUTC7 ( pull_down120 )
     ,.P140DIN ( P140DIN ) ,.P141DIN ( P141DIN ) ,.P146DIN ( P146DIN )
     ,.P147DIN ( P147DIN ) ,.P140ENO ( P140ENO ) ,.P141ENO ( P141ENO )
     ,.P146ENO ( P146ENO ) ,.P147ENO ( P147ENO ) ,.P140PUON ( P140PUON )
     ,.P141PUON ( P141PUON ) ,.P146PUON ( P146PUON ) ,.P147PUON ( P147PUON )
     ,.P140DOUT ( P140DOUT ) ,.P141DOUT ( P141DOUT ) ,.P146DOUT ( P146DOUT )
     ,.P147DOUT ( P147DOUT ) ,.P140ENI ( P140ENI ) ,.P141ENI ( P141ENI )
     ,.P146ENI ( P146ENI ) ,.P147ENI ( P147ENI ) ,.PIO140 ( PIO140 ) ,.PIO141 ( PIO141 )
     ,.PIO146 ( PIO146 ) ,.PIO147 ( PIO147 ) ,.EXOR ( PORT14EXOR )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_2.0/_macro/_local/kx4_pior_mf3_v2.00/_library/100821/kx4_piorv2.hdl
  KX4_PIORV2 pior (
    .PIOR0 ( PIOR0 ) ,.PIOR1 ( PIOR1 ) ,.PIOR2 ( PIOR2 ) ,.PIOR3 ( PIOR3 )
     ,.PIOR4 ( PIOR4 ) ,.TOUT00 ( TOUT00 ) ,.TOUT02 ( TOUT02 ) ,.TOUT03 ( TOUT03 )
     ,.TOUT04 ( TOUT04 ) ,.TOUT05 ( TOUT05 ) ,.TOUT06 ( TOUT06 ) ,.TOUT07 ( TOUT07 )
     ,.SOUT000 ( SOUT000 ) ,.SOUT002 ( SOUT002 ) ,.SOUT100 ( SOUT100 )
     ,.SOUT003 ( SOUT003 ) ,.SOUT013 ( SOUT013DLY ) ,.SCKO00 ( SCKO00 )
     ,.SCLO0 ( SCLO0 ) ,.SDAO0 ( SDAO0 ) ,.PCLBUZ0 ( PCLBUZ0 ) ,.PCLBUZ1 ( PCLBUZ1 )
     ,.P00EXINA ( P00EXINA ) ,.P01EXINA ( P01EXINA ) ,.P02EXINA ( P02EXINA )
     ,.P10EXINA ( P10EXINA ) ,.P03EXINA ( P03EXINA ) ,.P11EXINA ( P11EXINA )
     ,.P05EXINA ( P05EXINA ) ,.P13EXINA ( P13EXINA ) ,.P06EXINA ( P06EXINA )
     ,.P14EXINA ( P14EXINA ) ,.P12EXINA ( P12EXINA ) ,.P15EXINA ( P15EXINA )
     ,.P31EXINA ( P31EXINA ) ,.P16EXINA ( P16EXINA ) ,.P17EXINA ( P17EXINA )
     ,.P41EXINA ( P41EXINA ) ,.P42EXINA ( P42EXINA ) ,.P50EXINA ( P50EXINA )
     ,.P52EXINA ( P52EXINA ) ,.P60EXINA ( P60EXINA ) ,.P53EXINA ( P53EXINA )
     ,.P61EXINA ( P61EXINA ) ,.P55EXINA ( P55EXINA ) ,.P76EXINA ( P76EXINA )
     ,.P77EXINA ( P77EXINA ) ,.SEL64P ( SEL64P ) ,.SEL48P ( SEL48P ) ,.SEL52P ( SEL52P )
     ,.SEL44P ( SEL44P ) ,.SEL36P ( SEL36P ) ,.SEL40P ( SEL40P ) ,.SEL32P ( SEL32P )
     ,.SEL24P ( SEL24P ) ,.SEL38P ( SEL38P ) ,.SCKI00 ( SCKI00 ) ,.SEL30P ( SEL30P )
     ,.SEL20P ( SEL20P ) ,.TIN00 ( TIN00 ) ,.TIN02 ( TIN02 ) ,.TIN03 ( TIN03 )
     ,.TIN04 ( TIN04 ) ,.TIN05 ( TIN05 ) ,.TIN06 ( TIN06 ) ,.TIN07 ( TIN07 )
     ,.SIN00 ( SIN00 ) ,.SIN02 ( SIN02 ) ,.SIN10 ( SIN10 ) ,.SIN03 ( SIN03 )
     ,.INTP5EG ( INTP5EG ) ,.INTP10EG ( INTP10EG ) ,.INTP11EG ( INTP11EG )
     ,.SCLI0 ( SCLI0 ) ,.SDAI0 ( SDAI0 ) ,.P00EXOUTA ( P00EXOUTA ) ,.P01EXOUTB ( P01EXOUTB )
     ,.P02EXOUTA ( P02EXOUTA ) ,.P10EXOUTA ( P10EXOUTA ) ,.P03EXOUTB ( P03EXOUTB )
     ,.P11EXOUTB ( P11EXOUTB ) ,.P05EXOUTB ( P05EXOUTB ) ,.P13EXOUTB ( P13EXOUTB )
     ,.P06EXOUTB ( P06EXOUTB ) ,.P14EXOUTB ( P14EXOUTB ) ,.P10EXOUTB ( P10EXOUTB )
     ,.TXSAU ( TXSAU ) ,.P12EXOUTB ( P12EXOUTB ) ,.P13EXOUTA ( P13EXOUTA )
     ,.P13EXOUTC ( P13EXOUTC ) ,.P14EXOUTC ( P14EXOUTC ) ,.P15EXOUTB ( P15EXOUTB )
     ,.P31EXOUTB ( P31EXOUTB ) ,.P15EXOUTC ( P15EXOUTC ) ,.P31EXOUTC ( P31EXOUTC )
     ,.P16EXOUTA ( P16EXOUTA ) ,.P17EXOUTA ( P17EXOUTA ) ,.P17EXOUTB ( P17EXOUTB )
     ,.P41EXOUTB ( P41EXOUTB ) ,.P42EXOUTB ( P42EXOUTB ) ,.P51EXOUTA ( P51EXOUTA )
     ,.P55EXOUTA ( P55EXOUTA ) ,.P55EXOUTB ( P55EXOUTB ) ,.P60EXOUTB ( P60EXOUTB )
     ,.P61EXOUTB ( P61EXOUTB ) ,.P77EXOUTA ( P77EXOUTA ) ,.P140EXOUTB ( P140EXOUTB )
     ,.P141EXOUTB ( P141EXOUTB ) ,.BBSWPICA ( BBSWPICA ) ,.P10EXINB ( P10EXINB )
     ,.P10EXOUTC ( P10EXOUTC ) ,.P11EXOUTC ( P11EXOUTC )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/_ice/_macro/_eva/_kx4/_061/qlk0radaa32v1_eva.v
  QLK0RADAA32V1 adctl (
    .PCLK ( PCLKADC ) ,.PCLKRW ( PCLKRW ) ,.PRESETZ ( PRESADCZ ) ,.SCANCLK ( SCANCLK )
     ,.PADDR2 ( PADDR2 ) ,.PADDR1 ( PADDR1 ) ,.PADDR0 ( PADDR0 ) ,.PSEL1 ( PSELAD1 )
     ,.PSEL2 ( PSELAD2 ) ,.PWRITE ( PWRITE ) ,.PENABLE ( PENABLE ) ,.PWDATA15 ( MDW15 )
     ,.PWDATA14 ( MDW14 ) ,.PWDATA13 ( MDW13 ) ,.PWDATA12 ( MDW12 ) ,.PWDATA11 ( MDW11 )
     ,.PWDATA10 ( MDW10 ) ,.PWDATA9 ( MDW9 ) ,.PWDATA8 ( MDW8 ) ,.PWDATA7 ( MDW7 )
     ,.PWDATA6 ( MDW6 ) ,.PWDATA5 ( MDW5 ) ,.PWDATA4 ( MDW4 ) ,.PWDATA3 ( MDW3 )
     ,.PWDATA2 ( MDW2 ) ,.PWDATA1 ( MDW1 ) ,.PWDATA0 ( MDW0 ) ,.TTRG0 ( INTTM01 )
     ,.TTRG1 ( ADTRIG0 ) ,.TTRG2 ( TTRG2 ) ,.TTRG3 ( INTRTCI ) ,.ADEOCB ( ADEOCB )
     ,.ADSAR9 ( ADSAR9 ) ,.ADSAR8 ( ADSAR8 ) ,.ADSAR7 ( ADSAR7 ) ,.ADSAR6 ( ADSAR6 )
     ,.ADSAR5 ( ADSAR5 ) ,.ADSAR4 ( ADSAR4 ) ,.ADSAR3 ( ADSAR3 ) ,.ADSAR2 ( ADSAR2 )
     ,.ADSAR1 ( ADSAR1 ) ,.ADSAR0 ( ADSAR0 ) ,.SCANEN ( SCANEN ) ,.SCANMODE ( SCANMODE )
     ,.TESDBT ( TESDBT ) ,.REQPCLK ( REQPCLKAD ) ,.PRDATA15 ( PRDAD15 )
     ,.PRDATA14 ( PRDAD14 ) ,.PRDATA13 ( PRDAD13 ) ,.PRDATA12 ( PRDAD12 )
     ,.PRDATA11 ( PRDAD11 ) ,.PRDATA10 ( PRDAD10 ) ,.PRDATA9 ( PRDAD9 )
     ,.PRDATA8 ( PRDAD8 ) ,.PRDATA7 ( PRDAD7 ) ,.PRDATA6 ( PRDAD6 ) ,.PRDATA5 ( PRDAD5 )
     ,.PRDATA4 ( PRDAD4 ) ,.PRDATA3 ( PRDAD3 ) ,.PRDATA2 ( PRDAD2 ) ,.PRDATA1 ( PRDAD1 )
     ,.PRDATA0 ( PRDAD0 ) ,.INTAD ( INTAD ) ,.ADCLK ( ADCLK ) ,.ADPDB ( ADPDB )
     ,.ADCHSEL4 ( ADCHSEL4 ) ,.ADCHSEL3 ( ADCHSEL3 ) ,.ADCHSEL2 ( ADCHSEL2 )
     ,.ADCHSEL1 ( ADCHSEL1 ) ,.ADCHSEL0 ( ADCHSEL0 ) ,.ADBIONB ( ADBIONB )
     ,.ADS1 ( ADS1 ) ,.ADOFC ( ADOFC ) ,.ADCMP ( ADCMP ) ,.ADCPON ( ADCPON )
     ,.BG2ADEN ( BG2ADEN ) ,.BG2ADSEL ( BG2ADSEL ) ,.ADVSELMOD0 ( ADVSELMOD0 )
     ,.ADVSELMOD1 ( ADVSELMOD1 ) ,.ADGSELMOD ( ADGSELMOD ) ,.ADTESMOD0 ( ADTESMOD0 )
     ,.ADTESMOD1 ( ADTESMOD1 ) ,.ADTESMOD2 ( ADTESMOD2 ) ,.reg_adtyp ( reg_adtyp )
    
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_2.0/_macro/_local/_kx4_cap/kx4_capckgate_mf3_v1.00/_library/100927/kx4_capckgate.hdl
  KX4_CAPCKGATE capckgate (
    .BBMOSC ( BBMOSC ) ,.OSCOUTM ( OSCOUTM ) ,.BBHIOSC ( BBHIOSC ) ,.R32MOUT ( R32MOUT )
     ,.BBFMAIN ( BBFMAIN ) ,.FMAIN ( FMAIN ) ,.BBFSUB ( BBFSUB ) ,.FSUB ( FSUB )
     ,.BBFCLK ( BBFCLK ) ,.FCLKRT ( FCLKRT ) ,.BBFIL ( BBFIL ) ,.R15KOUT ( R15KOUT )
     ,.BBMODE ( BBMODE ) ,.SCANMODE ( SCANMODE )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_2.0/_macro/_local/_kx4_cap/kx4_capmux4_mf3_v1.00/_library/100826_noRAMext/kx4_capmux4.v
  KX4_CAPMUX4 capmux (
    .TTRG2 ( TTRG2 ) ,.INTRTC ( INTRTC ) ,.INTRTDISL ( INTRTDISL ) ,.INTRTDISR ( INTRTDISR )
     ,.BBCLKR ( BBCLKR ) ,.BBCLKM ( BBCLKM ) ,.BBREQPCLK ( BBREQPCLK )
     ,.BBCKSELR ( BBCKSELR ) ,.BBPRDATA15 ( BBPRDATA15 ) ,.BBPRDATA14 ( BBPRDATA14 )
     ,.BBPRDATA13 ( BBPRDATA13 ) ,.BBPRDATA12 ( BBPRDATA12 ) ,.BBPRDATA11 ( BBPRDATA11 )
     ,.BBPRDATA10 ( BBPRDATA10 ) ,.BBPRDATA9 ( BBPRDATA9 ) ,.BBPRDATA8 ( BBPRDATA8 )
     ,.BBPRDATA7 ( BBPRDATA7 ) ,.BBPRDATA6 ( BBPRDATA6 ) ,.BBPRDATA5 ( BBPRDATA5 )
     ,.BBPRDATA4 ( BBPRDATA4 ) ,.BBPRDATA3 ( BBPRDATA3 ) ,.BBPRDATA2 ( BBPRDATA2 )
     ,.BBPRDATA1 ( BBPRDATA1 ) ,.BBPRDATA0 ( BBPRDATA0 ) ,.BBWAITMEM ( BBWAITMEM )
     ,.BBWAIT56 ( BBWAIT56 ) ,.BBINT0 ( BBINT0 ) ,.BBINT1 ( BBINT1 ) ,.BBINT2 ( BBINT2 )
     ,.BBINT3 ( BBINT3 ) ,.BBINT4 ( BBINT4 ) ,.BBINT5 ( BBINT5 ) ,.BBINT6 ( BBINT6 )
     ,.BBINT7 ( BBINT7 ) ,.BBINT8 ( BBINT8 ) ,.BBINT9 ( BBINT9 ) ,.BBINT10 ( BBINT10 )
     ,.BBINT11 ( BBINT11 ) ,.BBINT12 ( BBINT12 ) ,.BBINT13 ( BBINT13 )
     ,.BBMODE ( BBMODE ) ,.BBSCANOUT ( BBSCANOUT ) ,.ADTRIG0 ( ADTRIG0 )
     ,.FRQ4EN ( FRQ4EN ) ,.BBCKSELM ( BBCKSELM ) ,.BBHIOON ( BBHIOON )
     ,.BBREGCTL ( BBREGCTL ) ,.BBCLKRL ( BBCLKRL ) ,.BBCLKRR ( BBCLKRR )
     ,.BBCLKML ( BBCLKML ) ,.BBCLKMR ( BBCLKMR ) ,.BBREQPCLKL ( BBREQPCLKL )
     ,.BBREQPCLKR ( BBREQPCLKR ) ,.BBCKSELRL ( BBCKSELRL ) ,.BBCKSELRR ( BBCKSELRR )
     ,.BBPRDATA15L ( BBPRDATA15L ) ,.BBPRDATA12R ( BBPRDATA12R ) ,.BBPRDATA15R ( BBPRDATA15R )
     ,.BBPRDATA14L ( BBPRDATA14L ) ,.BBPRDATA11R ( BBPRDATA11R ) ,.BBPRDATA14R ( BBPRDATA14R )
     ,.BBPRDATA13L ( BBPRDATA13L ) ,.BBPRDATA10R ( BBPRDATA10R ) ,.BBPRDATA13R ( BBPRDATA13R )
     ,.BBPRDATA12L ( BBPRDATA12L ) ,.BBPRDATA11L ( BBPRDATA11L ) ,.BBPRDATA10L ( BBPRDATA10L )
     ,.BBPRDATA9L ( BBPRDATA9L ) ,.BBPRDATA6R ( BBPRDATA6R ) ,.BBPRDATA9R ( BBPRDATA9R )
     ,.BBPRDATA8L ( BBPRDATA8L ) ,.BBPRDATA5R ( BBPRDATA5R ) ,.BBPRDATA8R ( BBPRDATA8R )
     ,.BBPRDATA7L ( BBPRDATA7L ) ,.BBPRDATA4R ( BBPRDATA4R ) ,.BBPRDATA7R ( BBPRDATA7R )
     ,.BBPRDATA6L ( BBPRDATA6L ) ,.BBPRDATA3R ( BBPRDATA3R ) ,.BBPRDATA5L ( BBPRDATA5L )
     ,.BBPRDATA2R ( BBPRDATA2R ) ,.BBPRDATA4L ( BBPRDATA4L ) ,.BBPRDATA1R ( BBPRDATA1R )
     ,.BBPRDATA3L ( BBPRDATA3L ) ,.BBPRDATA0R ( BBPRDATA0R ) ,.BBPRDATA2L ( BBPRDATA2L )
     ,.BBPRDATA1L ( BBPRDATA1L ) ,.BBPRDATA0L ( BBPRDATA0L ) ,.BBWAITMEML ( BBWAITMEML )
     ,.BBWAITMEMR ( BBWAITMEMR ) ,.BBWAIT56L ( BBWAIT56L ) ,.BBWAIT56R ( BBWAIT56R )
     ,.BBINT0L ( BBINT0L ) ,.BBINT0R ( BBINT0R ) ,.BBINT3L ( BBINT3L )
     ,.BBINT1L ( BBINT1L ) ,.BBINT1R ( BBINT1R ) ,.BBINT4L ( BBINT4L )
     ,.BBINT2L ( BBINT2L ) ,.BBINT2R ( BBINT2R ) ,.BBINT5L ( BBINT5L )
     ,.BBINT3R ( BBINT3R ) ,.BBINT6L ( BBINT6L ) ,.BBINT4R ( BBINT4R )
     ,.BBINT7L ( BBINT7L ) ,.BBINT5R ( BBINT5R ) ,.BBINT8L ( BBINT8L )
     ,.BBINT6R ( BBINT6R ) ,.BBINT9L ( BBINT9L ) ,.BBINT7R ( BBINT7R )
     ,.BBINT8R ( BBINT8R ) ,.BBINT9R ( BBINT9R ) ,.BBINT10L ( BBINT10L )
     ,.BBINT10R ( BBINT10R ) ,.BBINT13L ( BBINT13L ) ,.BBINT11L ( BBINT11L )
     ,.BBINT11R ( BBINT11R ) ,.BBINT12L ( BBINT12L ) ,.BBINT12R ( BBINT12R )
     ,.BBINT13R ( BBINT13R ) ,.BBMODEL ( BBMODEL ) ,.BBMODER ( BBMODER )
     ,.BBSCANOUTL ( BBSCANOUTL ) ,.BBSCANOUTR ( BBSCANOUTR ) ,.ADTRIG0L ( ADTRIG0L )
     ,.ADTRIG0R ( ADTRIG0R ) ,.ADTRIG1L ( ADTRIG1L ) ,.ADTRIG1R ( ADTRIG1R )
     ,.FRQ4ENL ( FRQ4ENL ) ,.FRQ4ENR ( FRQ4ENR ) ,.BBCKSELML ( BBCKSELML )
     ,.BBCKSELMR ( BBCKSELMR ) ,.BBHIOONL ( BBHIOONL ) ,.BBHIOONR ( BBHIOONR )
     ,.BBREGCTLL ( BBREGCTLL ) ,.BBREGCTLR ( BBREGCTLR )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_2.0/_macro/_local/_kx4_cap/kx4_caplrio_mf3_v1.00/_library/100904/kx4_caplio.v_RAMext
  KX4_CAPLIO capl (
    .SELIN1B5V ( P40SELIN1B5V ) ,.BBMOSC ( BBMOSC ) ,.BBHIOSC ( BBHIOSC )
     ,.BBFMAIN ( BBFMAIN ) ,.BBFSUB ( BBFSUB ) ,.BBFCLK ( BBFCLK ) ,.BBFIL ( BBFIL )
     ,.BBCLKRIL ( BBCLKRL ) ,.BBCLKMIL ( BBCLKML ) ,.SYSRESB ( SYSRESB )
     ,.RESETB ( RESETB ) ,.RESB ( RESB ) ,.STPBCKBT ( STPBCKBT ) ,.RSTS ( RSTS )
     ,.RESSTP ( RESSTP ) ,.FMXST ( FMXST ) ,.SUBCKST ( SUBCKST ) ,.BCKHSEN ( BCKHSEN )
     ,.BBCKSTR ( BBCKSTR ) ,.BBCKSTM ( BBCKSTM ) ,.BBPWRITE ( BBPWRITE )
     ,.BBPENABLE ( BBPENABLE ) ,.BBMA10 ( BBMA10 ) ,.BBMA9 ( BBMA9 ) ,.BBMA8 ( BBMA8 )
     ,.BBMA7 ( BBMA7 ) ,.BBMA6 ( BBMA6 ) ,.BBMA5 ( BBMA5 ) ,.BBMA4 ( BBMA4 )
     ,.BBMA3 ( BBMA3 ) ,.BBMA2 ( BBMA2 ) ,.BBMA1 ( BBMA1 ) ,.BBMA0 ( BBMA0 )
     ,.MDWFLRO15 ( MDWFLRO15 ) ,.MDWFLRO14 ( MDWFLRO14 ) ,.MDWFLRO13 ( MDWFLRO13 )
     ,.MDWFLRO12 ( MDWFLRO12 ) ,.MDWFLRO11 ( MDWFLRO11 ) ,.MDWFLRO10 ( MDWFLRO10 )
     ,.MDWFLRO9 ( MDWFLRO9 ) ,.MDWFLRO8 ( MDWFLRO8 ) ,.MDWFLRO7 ( MDWFLRO7 )
     ,.MDWFLRO6 ( MDWFLRO6 ) ,.MDWFLRO5 ( MDWFLRO5 ) ,.MDWFLRO4 ( MDWFLRO4 )
     ,.MDWFLRO3 ( MDWFLRO3 ) ,.MDWFLRO2 ( MDWFLRO2 ) ,.MDWFLRO1 ( MDWFLRO1 )
     ,.MDWFLRO0 ( MDWFLRO0 ) ,.BBNVM1 ( BBNVM1 ) ,.BBNVM2 ( BBNVM2 ) ,.SVSTOP ( SVSTOP )
     ,.SVPERI0 ( SVPERI0 ) ,.SVPERI1 ( SVPERI1 ) ,.SCANMODE ( SCANMODE )
     ,.SCANEN ( SCANEN ) ,.SCANIN ( SCANIN ) ,.BBTESSCAN1 ( TESSCAN1 )
     ,.BBTESINST ( BBTESINST ) ,.OPTIDDQ ( OPTIDDQ ) ,.OPTEXCCK ( OPTEXCCK )
     ,.TESDBT2 ( TESDBT2 ) ,.TESDBT ( TESDBT ) ,.SEL08P ( SEL08P ) ,.SLMEM ( SLMEM )
     ,.FCHRAM ( FCHRAM ) ,.WDOP ( WDOP ) ,.BBSTN ( STN ) ,.MODE0 ( MODE0 )
     ,.MODE1 ( MODE1 ) ,.GDRAMWR ( GDRAMWR ) ,.BBMA15 ( BBMA15 ) ,.BBMA14 ( BBMA14 )
     ,.BBMA13 ( BBMA13 ) ,.BBMA12 ( BBMA12 ) ,.BBMA11 ( BBMA11 ) ,.BBRPERRIL ( BBRPERR )
     ,.BBREQPCLKIL ( BBREQPCLKL ) ,.BBCKSELRIL ( BBCKSELRL ) ,.BBPRDATA15IL ( BBPRDATA15L )
     ,.BBPRDATA14IL ( BBPRDATA14L ) ,.BBPRDATA13IL ( BBPRDATA13L ) ,.BBPRDATA12IL ( BBPRDATA12L )
     ,.BBPRDATA11IL ( BBPRDATA11L ) ,.BBPRDATA10IL ( BBPRDATA10L ) ,.BBPRDATA9IL ( BBPRDATA9L )
     ,.BBPRDATA8IL ( BBPRDATA8L ) ,.BBPRDATA7IL ( BBPRDATA7L ) ,.BBPRDATA6IL ( BBPRDATA6L )
     ,.BBPRDATA5IL ( BBPRDATA5L ) ,.BBPRDATA4IL ( BBPRDATA4L ) ,.BBPRDATA3IL ( BBPRDATA3L )
     ,.BBPRDATA2IL ( BBPRDATA2L ) ,.BBPRDATA1IL ( BBPRDATA1L ) ,.BBPRDATA0IL ( BBPRDATA0L )
     ,.BBWAITMEMIL ( BBWAITMEML ) ,.BBWAIT56IL ( BBWAIT56L ) ,.BBINT0IL ( BBINT0L )
     ,.BBINT1IL ( BBINT1L ) ,.BBINT2IL ( BBINT2L ) ,.BBINT3IL ( BBINT3L )
     ,.BBINT4IL ( BBINT4L ) ,.BBINT5IL ( BBINT5L ) ,.BBINT6IL ( BBINT6L )
     ,.BBINT7IL ( BBINT7L ) ,.BBINT8IL ( BBINT8L ) ,.BBINT9IL ( BBINT9L )
     ,.BBINT10IL ( BBINT10L ) ,.BBINT11IL ( BBINT11L ) ,.BBINT12IL ( BBINT12L )
     ,.BBINT13IL ( BBINT13L ) ,.BBMODEIL ( BBMODEL ) ,.BBSCANOUTIL ( BBSCANOUTL )
     ,.ADTRIG0IL ( ADTRIG0L ) ,.ADTRIG1IL ( ADTRIG1L ) ,.FRQ4ENIL ( FRQ4ENL )
     ,.INTRTDISIL ( INTRTDISL ) ,.BBCKSELMIL ( BBCKSELML ) ,.BBHIOONIL ( BBHIOONL )
     ,.BBREGCTLIL ( BBREGCTLL )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_2.0/_macro/_local/_kx4_cap/kx4_caplrio_mf3_v1.00/_library/101109/kx4_caprio.v_noRAMext
  KX4_CAPRIO capr (
    .SELIN1B5V ( P147SELIN1B5V ) ,.SCANCLK ( SCANCLK ) ,.BBMOSC ( BBMOSC )
     ,.BBHIOSC ( BBHIOSC ) ,.BBFMAIN ( BBFMAIN ) ,.BBFSUB ( BBFSUB ) ,.BBFCLK ( BBFCLK )
     ,.BBFIL ( BBFIL ) ,.BBCLKRIR ( BBCLKRR ) ,.BBCLKMIR ( BBCLKMR ) ,.SYSRESB ( SYSRESB )
     ,.RESETB ( RESETB ) ,.RESB ( RESB ) ,.STPBCKBT ( STPBCKBT ) ,.RSTS ( RSTS )
     ,.RESSTP ( RESSTP ) ,.FMXST ( FMXST ) ,.SUBCKST ( SUBCKST ) ,.BCKHSEN ( BCKHSEN )
     ,.BBCKSTR ( BBCKSTR ) ,.BBCKSTM ( BBCKSTM ) ,.BBPWRITE ( BBPWRITE )
     ,.BBPENABLE ( BBPENABLE ) ,.BBMA10 ( BBMA10 ) ,.BBMA9 ( BBMA9 ) ,.BBMA8 ( BBMA8 )
     ,.BBMA7 ( BBMA7 ) ,.BBMA6 ( BBMA6 ) ,.BBMA5 ( BBMA5 ) ,.BBMA4 ( BBMA4 )
     ,.BBMA3 ( BBMA3 ) ,.BBMA2 ( BBMA2 ) ,.BBMA1 ( BBMA1 ) ,.BBMA0 ( BBMA0 )
     ,.MDWFLRO15 ( MDWFLRO15 ) ,.MDWFLRO14 ( MDWFLRO14 ) ,.MDWFLRO13 ( MDWFLRO13 )
     ,.MDWFLRO12 ( MDWFLRO12 ) ,.MDWFLRO11 ( MDWFLRO11 ) ,.MDWFLRO10 ( MDWFLRO10 )
     ,.MDWFLRO9 ( MDWFLRO9 ) ,.MDWFLRO8 ( MDWFLRO8 ) ,.MDWFLRO7 ( MDWFLRO7 )
     ,.MDWFLRO6 ( MDWFLRO6 ) ,.MDWFLRO5 ( MDWFLRO5 ) ,.MDWFLRO4 ( MDWFLRO4 )
     ,.MDWFLRO3 ( MDWFLRO3 ) ,.MDWFLRO2 ( MDWFLRO2 ) ,.MDWFLRO1 ( MDWFLRO1 )
     ,.MDWFLRO0 ( MDWFLRO0 ) ,.BBNVM1 ( BBNVM1 ) ,.BBNVM2 ( BBNVM2 ) ,.SVSTOP ( SVSTOP )
     ,.SVPERI0 ( SVPERI0 ) ,.SVPERI1 ( SVPERI1 ) ,.SCANMODE ( SCANMODE )
     ,.SCANEN ( SCANEN ) ,.SCANIN ( SCANIN ) ,.BBTESSCAN1 ( TESSCAN1 )
     ,.BBTESINST ( BBTESINST ) ,.OPTIDDQ ( OPTIDDQ ) ,.OPTEXCCK ( OPTEXCCK )
     ,.TESDBT2 ( TESDBT2 ) ,.TESDBT ( TESDBT ) ,.SEL08P ( SEL08P ) ,.BBSELSFR1 ( BBSELSFR1 )
     ,.BBSELSFR2 ( BBSELSFR2 ) ,.BBEXIP12 ( P12EXINB ) ,.BBEXIP10 ( P10EXINB )
     ,.BBEXIP11 ( P11EXINA ) ,.BBREQPCLKIR ( BBREQPCLKR ) ,.BBCKSELRIR ( BBCKSELRR )
     ,.BBPRDATA15IR ( BBPRDATA15R ) ,.BBPRDATA14IR ( BBPRDATA14R ) ,.BBPRDATA13IR ( BBPRDATA13R )
     ,.BBPRDATA12IR ( BBPRDATA12R ) ,.BBPRDATA11IR ( BBPRDATA11R ) ,.BBPRDATA10IR ( BBPRDATA10R )
     ,.BBPRDATA9IR ( BBPRDATA9R ) ,.BBPRDATA8IR ( BBPRDATA8R ) ,.BBPRDATA7IR ( BBPRDATA7R )
     ,.BBPRDATA6IR ( BBPRDATA6R ) ,.BBPRDATA5IR ( BBPRDATA5R ) ,.BBPRDATA4IR ( BBPRDATA4R )
     ,.BBPRDATA3IR ( BBPRDATA3R ) ,.BBPRDATA2IR ( BBPRDATA2R ) ,.BBPRDATA1IR ( BBPRDATA1R )
     ,.BBPRDATA0IR ( BBPRDATA0R ) ,.BBWAITMEMIR ( BBWAITMEMR ) ,.BBWAIT56IR ( BBWAIT56R )
     ,.BBINT0IR ( BBINT0R ) ,.BBINT1IR ( BBINT1R ) ,.BBINT2IR ( BBINT2R )
     ,.BBINT3IR ( BBINT3R ) ,.BBINT4IR ( BBINT4R ) ,.BBINT5IR ( BBINT5R )
     ,.BBINT6IR ( BBINT6R ) ,.BBINT7IR ( BBINT7R ) ,.BBINT8IR ( BBINT8R )
     ,.BBINT9IR ( BBINT9R ) ,.BBINT10IR ( BBINT10R ) ,.BBINT11IR ( BBINT11R )
     ,.BBINT12IR ( BBINT12R ) ,.BBINT13IR ( BBINT13R ) ,.BBMODEIR ( BBMODER )
     ,.BBSCANOUTIR ( BBSCANOUTR ) ,.ADTRIG0IR ( ADTRIG0R ) ,.ADTRIG1IR ( ADTRIG1R )
     ,.FRQ4ENIR ( FRQ4ENR ) ,.INTRTDISIR ( INTRTDISR ) ,.BBCKSELMIR ( BBCKSELMR )
     ,.BBHIOONIR ( BBHIOONR ) ,.BBREGCTLIR ( BBREGCTLR ) ,.BBEXAD10 ( BBEXAD10 )
     ,.BBEXAD11 ( BBEXAD11 ) ,.BBEXAD12 ( BBEXAD12 ) ,.BBEXOR10 ( BBEXOR10 )
     ,.BBEXOR11 ( BBEXOR11 ) ,.BBEXOR12 ( BBEXOR12 ) ,.BBSFDIS1 ( BBSFDIS1 )
     ,.BBSWPPT1 ( BBSWPPT1 ) ,.BBSWPICA ( BBSWPICA ) ,.BBISC ( BBISC )
    
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/HMG_IOBUF_SS3_KX4V2_mf3_v2.00_LR4.2.16_20100924/_misc/lib/MF3/cmos1_2.1V/verilog/QICAP035H5H.v
  QICAP035H5H capadl (
    .ADINLBB5V ( ADINLBB5V )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/HMG_IOBUF_SS3_KX4V2_mf3_v2.00_LR4.2.16_20100924/_misc/lib/MF3/cmos1_2.1V/verilog/QICAP025H5H.v
  QICAP025H5H capadr (
    .ADINLBB5V ( ADINL5V )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/tbfilter1x2_mf3_v1.02_20100730/_misc/lib/MF3/cmos1_2.1V/verilog/TBFILTER1X2.v
  TBFILTER1X2 dmydly50n (
    .N01 ( DLY50NO ) ,.H01 ( P13EXINA )
  ) ;
  // Refer to /proj/78k0r_11/78k0r_kx4/top_1.0/_macro/_hard/qahnfi4bn300nv1_mf3_v1.11/_misc/lib/MF3/cmos1_2.1V/verilog/QAHNFI4BN300NV1.v
  QAHNFI4BN300NV1 dmydly300n (
    .NFOUT ( DLY300NO ) ,.NFIN ( P14EXINA )
  ) ;
  // Refer to /proj/78k0r_16/ss3rd/_macro/_1_local_release/_hard/HMG_IOBUF_SS3_KX4V2_mf3_v2.00_LR4.2.16_20100924/_misc/lib/MF3/cmos1_2.1V/verilog/QAHRES0CV1.v
  QAHRES0CV1 vppts1_res (
    .VPPTSIN ( VPPTS1 ) ,.VPPTSOUT ( VPPTS1_CP )
  ) ;
endmodule
/********************************************************************************/
/* K0R CPUEVA Macro                                                           	*/
/*                                      Made K.Ishihara K.tanaka K.kawai        */
/********************************************************************************/
/* Ver1.00  New                                                                 */
/* Ver1.50  Add FLREAD                                2007.05.30 K.Tanaka       */
/*              FCHRAM                                2007.05.30 K.Tanaka       */
/*              mem_access                            2007.05.30 K.Tanaka       */
/*              stbst                                 2007.07.02 K.Tanaka       */
/* Ver1.51  Add OCDMOD                                2007.11.30 K.Tanaka       */
/* Ver1.52  Modified MONMD Signal during svmod        2008.02.26 K.Tanaka       */
/* Ver2.00  ��������̸�ľ��                        2008.01.16 K.Ishihara	*/
/*            ADR:���ɥ쥹�黻���adrout_pc,adrout_ma,adrout_sub�ˣ�ʬ��	*/
/*������������ADR:SLFLASH���Ϥη�ϩ���®��					*/
/*������������ADR:imdr�����Ϸ�ϩ�򺬸��ǥޥ���					*/
/*������������ADR:����������ϩ��intclk_on�ο���ǥ����ƥ���			*/
/*������������ALU:ALU��5ʬ�䡢exeout,muluout,transout,transin,bitshout		*/
/*������������ALU:imdr,���ѥ쥸�����������Ϸ�ϩ�򺬸��ǥޥ���			*/
/* Ver2.01  Modified CPUMISAL Signal                  2008.08.29 K.Tanaka       */
/* Ver3.00  ����ή��ϩ���(Ver2.00�ɲ�ʬ)					*/
/*	    DataFlash�����������Υ������ȵ�ǽ�ɲ�				*/
/*	    ������ȯ������ʬ�����ѹ�						*/
/*	    ���ɥ쥹�Х��Υ����ƥ��󥰲�ϩ�ɲ�					*/
/*      2010.01.21                                                              */
/*              DataFlash�����������DMAž����ޥ���                            */
/*              - dmaack��������sldfwait_pre�ɲ�                                */
/*              PC�˥��եȥ֥쥤������ʬ�����ɲ�(BFA)                           */
/*              - softbrk_sub������ɲ�                                         */
/*      2010.01.26                                                              */
/*		PCʬ����ϩ��SVMOD�ˤ��ʬ�������ɲ�				*/
/*      2010.01.29                                                              */
/*		intack��WED�������ɲ�(���Ҥδ�ά��)				*/
/*      2010.02.02								*/
/* 		- OCDʬ����︫ľ��						*/
/*		  (monmd,ivack,softbrk_sub)->(monmd)				*/
/*		  softbrk_sub�������						*/
/*      2010.02.03								*/
/*		- CRC�黻��(modectl)�����HALT���������ɲ�(CRCHLTEN)		*/
/*      2010.02.04								*/
/*		- DataFlash�꡼�ɥ����ߥ󥰿�����ѹ�				*/
/*      2010.02.05								*/
/*		- DFlash vs 2ndSFR �ζ����б�					*/
/*		  �ߤ��Υ������Ȥ�ȯ�������Ȥ������Υ������ȿ����ޥ�������	*/
/*      2010.02.06								*/
/*		- ADR���ؤ�WEDü�� WED/wed �����ߤ��Ƥ������� wed ������	*/
/*      2010.02.10								*/
/*		- intack��MONMD��ͭ���ˤʤ�褦�������ɲ�			*/
/*		- BASECK -> BASECKHS(�ޥ���TOP)					*/
/*		- imdr_groupA�򥳥��ȥ�����(��³�褬�ʤ�)			*/
/*		- cpu�꡼�ɥХ�����ɥ�����������RVEON���Х��˾��褦�˽���	*/
/********************************************************************************/
module QLK0RCPUEVA0V3(
	PC19, PC18, PC17, PC16, PC15, PC14, PC13, PC12, PC11, PC10, PC9, PC8, PC7, PC6, PC5, PC4, PC3, PC2, PC1, PC0,
	PA19, PA18, PA17, PA16, PA15, PA14, PA13, PA12, PA11, PA10, PA9, PA8, PA7, PA6, PA5, PA4, PA3, PA2,
	PID31, PID30, PID29, PID28, PID27, PID26, PID25, PID24, PID23, PID22, PID21, PID20, PID19, PID18, PID17, PID16,
	PID15, PID14, PID13, PID12, PID11, PID10, PID9, PID8, PID7, PID6, PID5, PID4, PID3, PID2, PID1, PID0,
	MA15, MA14, MA13, MA12, MA11, MA10, MA9, MA8, MA7, MA6, MA5, MA4, MA3, MA2, MA1, MA0,
	DMAMA15, DMAMA14, DMAMA13, DMAMA12, DMAMA11, DMAMA10, DMAMA9, DMAMA8, DMAMA7, DMAMA6, DMAMA5,
	DMAMA4, DMAMA3, DMAMA2, DMAMA1, DMAMA0, DMARQ, DMAACK, DMARD, DMAWR, DMAWDOP, DMAEN,
	SLMEM, SLFLASH, SLEXM, SLBMEM, SLIRAM, HLTST, STPST, STBEN,
	MDR15, MDR14, MDR13, MDR12, MDR11, MDR10, MDR9, MDR8, MDR7, MDR6, MDR5, MDR4, MDR3, MDR2, MDR1, MDR0,
	MDW15, MDW14, MDW13, MDW12, MDW11, MDW10, MDW9, MDW8, MDW7, MDW6, MDW5, MDW4, MDW3, MDW2, MDW1, MDW0,
	BITEN7, BITEN6, BITEN5, BITEN4, BITEN3, BITEN2, BITEN1, BITEN0,
	CPUWR, CPURD, WDOP, WDWR, EXMA3, EXMA2, EXMA1, EXMA0,
	VCOUT6, VCOUT5, VCOUT4, VCOUT3, VCOUT2, VCOUT1,
	INTDBG, INTNMI, INTRQ3, INTRQ2, INTRQ1, INTRQ0, INTACK, SKIPEXE, MONMD, MONMDSTP, SOFTBRK, BRKMSK,
	WAITMEM, WAITFL, WAITMOD, WAITEXM, DMAWAIT, OCDWAIT,
	FLSIZE3, FLSIZE2, FLSIZE1, FLSIZE0, BFSIZE3, BFSIZE2, BFSIZE1, BFSIZE0,
	RAMSIZE7, RAMSIZE6, RAMSIZE5, RAMSIZE4, RAMSIZE3, RAMSIZE2, RAMSIZE1, RAMSIZE0,
	BMSIZE3, BMSIZE2, BMSIZE1, BMSIZE0,
	WAIT2ND7, WAIT2ND6, WAIT2ND5, WAIT2ND4, WAIT2ND3, WAIT2ND2, WAIT2ND1, WAIT2ND0,
	FLREAD, FCHRAM,
// for EVA
        WAITFL2, ICEWAITMEM,
        SVI, SVVCOUT7, SVVCOUT6, SVVCOUT5, SVVCOUT4, SVVCOUT3, SVVCOUT2, SVVCOUT1, SVVCOUT0,
        SVINTACK, SVMOD, SVMODF,
        ALT1, ALT2,
        SP15, SP14, SP13, SP12, SP11, SP10, SP9, SP8, SP7, SP6, SP5, SP4, SP3, SP2, SP1, SP0,
        SPINC, SPDEC, IDPOP,
        ICECSGREGU, ICECSGREGA, ICEIFA4, ICEIFA3, ICEIFA2,
        ICEDO31, ICEDO30, ICEDO29, ICEDO28, ICEDO27, ICEDO26, ICEDO25, ICEDO24,
        ICEDO23, ICEDO22, ICEDO21, ICEDO20, ICEDO19, ICEDO18, ICEDO17, ICEDO16,
        ICEDO15, ICEDO14, ICEDO13, ICEDO12, ICEDO11, ICEDO10, ICEDO9, ICEDO8,
        ICEDO7, ICEDO6, ICEDO5, ICEDO4, ICEDO3, ICEDO2, ICEDO1, ICEDO0,
        FLREADB3, FLREADB2, FLREADB1, FLREADB0,
        IMDR15, IMDR14, IMDR13, IMDR12, IMDR11, IMDR10, IMDR9, IMDR8,
        IMDR7, IMDR6, IMDR5, IMDR4, IMDR3, IMDR2, IMDR1, IMDR0,
        IDADR31, IDADR30, IDADR29, IDADR28, IDADR27, IDADR26, IDADR25, IDADR24,
        IDADR23, IDADR22, IDADR21, IDADR20, IDADR19, IDADR18, IDADR17, IDADR16,
        IDADR15, IDADR14, IDADR13, IDADR12, IDADR11, IDADR10, IDADR9, IDADR8,
        IDADR7, IDADR6, IDADR5, IDADR4, IDADR3, IDADR2, IDADR1, IDADR0,
        STAGEADR1, STAGEADR0,
        PREFIX, PCWAITF,
        ICEMSKNMI, ICEMSKDBG,
        CPUMASK, CPUMISAL, SPREL,
        // Ver1.51
        OCDMOD,
//
	PSELCPU, PSELBCD, CPUSTART, /*DECDYCUT,*/ BASECKHS, RESB, SCANMODE,
	DFSIZE1, DFSIZE0, DFLEN, SLDFLASH, DRDCLK,
	WED, FLSPM, GOFIRM,
	GATEAD1, GATEAD2, GATEAD3,
	MONPC19, MONPC18, MONPC17, MONPC16, MONPC15, MONPC14, MONPC13, MONPC12, MONPC11, MONPC10,
	MONPC9, MONPC8, MONPC7, MONPC6, MONPC5, MONPC4, MONPC3, MONPC2, MONPC1, MONPC0,
	MONMA15, MONMA14, MONMA13, MONMA12, MONMA11, MONMA10,
	MONMA9, MONMA8, MONMA7, MONMA6, MONMA5, MONMA4, MONMA3, MONMA2, MONMA1, MONMA0,
	MONMDR15, MONMDR14, MONMDR13, MONMDR12, MONMDR11, MONMDR10,
	MONMDR9, MONMDR8, MONMDR7, MONMDR6, MONMDR5, MONMDR4, MONMDR3, MONMDR2, MONMDR1, MONMDR0,
	MONMDW15, MONMDW14, MONMDW13, MONMDW12, MONMDW11, MONMDW10,
	MONMDW9, MONMDW8, MONMDW7, MONMDW6, MONMDW5, MONMDW4, MONMDW3, MONMDW2, MONMDW1, MONMDW0, 
	CRCHLTEN
	);

	output	PC19, PC18, PC17, PC16, PC15, PC14, PC13, PC12, PC11, PC10, PC9, PC8, PC7, PC6, PC5, PC4, PC3, PC2, PC1, PC0;
	output	PA19, PA18, PA17, PA16, PA15, PA14, PA13, PA12, PA11, PA10, PA9, PA8, PA7, PA6, PA5, PA4, PA3, PA2;
	output	MA15, MA14, MA13, MA12, MA11, MA10, MA9, MA8, MA7, MA6, MA5, MA4, MA3, MA2, MA1, MA0;
	output	DMAACK;
	output	SLMEM, SLFLASH, SLEXM, SLBMEM, SLIRAM;
	output	HLTST, STPST;
	output	STBEN;
	output	MDW15, MDW14, MDW13, MDW12, MDW11, MDW10, MDW9, MDW8, MDW7, MDW6, MDW5, MDW4, MDW3, MDW2, MDW1, MDW0;
	output	BITEN7, BITEN6, BITEN5, BITEN4, BITEN3, BITEN2, BITEN1, BITEN0;
	output	CPUWR, CPURD, WDOP, WDWR;
	output	EXMA3, EXMA2, EXMA1, EXMA0;
	output	INTACK;
	output	SKIPEXE;
	output	MONMD, MONMDSTP;
	output	SOFTBRK, BRKMSK;
	output	DMAWAIT, OCDWAIT;
	output	FLREAD, FCHRAM;
	output	SLDFLASH, DRDCLK;
	output	MONPC19, MONPC18, MONPC17, MONPC16, MONPC15, MONPC14, MONPC13, MONPC12, MONPC11, MONPC10;
	output	MONPC9, MONPC8, MONPC7, MONPC6, MONPC5, MONPC4, MONPC3, MONPC2, MONPC1, MONPC0;
	output	MONMA15, MONMA14, MONMA13, MONMA12, MONMA11, MONMA10;
	output	MONMA9, MONMA8, MONMA7, MONMA6, MONMA5, MONMA4, MONMA3, MONMA2, MONMA1, MONMA0;
	output	MONMDR15, MONMDR14, MONMDR13, MONMDR12, MONMDR11, MONMDR10;
	output	MONMDR9, MONMDR8, MONMDR7, MONMDR6, MONMDR5, MONMDR4, MONMDR3, MONMDR2, MONMDR1, MONMDR0;
	output	MONMDW15, MONMDW14, MONMDW13, MONMDW12, MONMDW11, MONMDW10;
	output	MONMDW9, MONMDW8, MONMDW7, MONMDW6, MONMDW5, MONMDW4, MONMDW3, MONMDW2, MONMDW1, MONMDW0;

// for EVA
        output  SVINTACK, SVMOD, SVMODF;
        output  ALT1, ALT2;
        output  SP15, SP14, SP13, SP12, SP11, SP10, SP9, SP8, SP7, SP6, SP5, SP4, SP3, SP2, SP1, SP0;
        output  SPINC, SPDEC, IDPOP;
        output  ICEDO31, ICEDO30, ICEDO29, ICEDO28, ICEDO27, ICEDO26, ICEDO25, ICEDO24;
        output  ICEDO23, ICEDO22, ICEDO21, ICEDO20, ICEDO19, ICEDO18, ICEDO17, ICEDO16;
        output  ICEDO15, ICEDO14, ICEDO13, ICEDO12, ICEDO11, ICEDO10, ICEDO9, ICEDO8;
        output  ICEDO7, ICEDO6, ICEDO5, ICEDO4, ICEDO3, ICEDO2, ICEDO1, ICEDO0;
        output  FLREADB3, FLREADB2, FLREADB1, FLREADB0;
        output  IMDR15, IMDR14, IMDR13, IMDR12, IMDR11, IMDR10, IMDR9, IMDR8;
        output  IMDR7, IMDR6, IMDR5, IMDR4, IMDR3, IMDR2, IMDR1, IMDR0;
        output  IDADR31, IDADR30, IDADR29, IDADR28, IDADR27, IDADR26, IDADR25, IDADR24;
        output  IDADR23, IDADR22, IDADR21, IDADR20, IDADR19, IDADR18, IDADR17, IDADR16;
        output  IDADR15, IDADR14, IDADR13, IDADR12, IDADR11, IDADR10, IDADR9, IDADR8;
        output  IDADR7, IDADR6, IDADR5, IDADR4, IDADR3, IDADR2, IDADR1, IDADR0;
        output  STAGEADR1, STAGEADR0;
        output  PREFIX, PCWAITF;
        output  CPUMASK, CPUMISAL, SPREL;
//

	input	PID31, PID30, PID29, PID28, PID27, PID26, PID25, PID24, PID23, PID22, PID21, PID20, PID19, PID18, PID17, PID16;
	input	PID15, PID14, PID13, PID12, PID11, PID10, PID9, PID8, PID7, PID6, PID5, PID4, PID3, PID2, PID1, PID0;
	input	DMAMA15, DMAMA14, DMAMA13, DMAMA12, DMAMA11, DMAMA10, DMAMA9, DMAMA8, DMAMA7, DMAMA6, DMAMA5;
	input	DMAMA4, DMAMA3, DMAMA2, DMAMA1, DMAMA0;
	input	DMARQ, DMARD, DMAWR, DMAWDOP, DMAEN;
	input	MDR15, MDR14, MDR13, MDR12, MDR11, MDR10, MDR9, MDR8, MDR7, MDR6, MDR5, MDR4, MDR3, MDR2, MDR1, MDR0;
	input	VCOUT6, VCOUT5, VCOUT4, VCOUT3, VCOUT2, VCOUT1;
	input	INTDBG, INTNMI, INTRQ3, INTRQ2, INTRQ1, INTRQ0;
	input	WAITMEM, WAITFL, WAITMOD, WAITEXM;
	input	FLSIZE3, FLSIZE2, FLSIZE1, FLSIZE0;
	input	BFSIZE3, BFSIZE2, BFSIZE1, BFSIZE0;
	input	RAMSIZE7, RAMSIZE6, RAMSIZE5, RAMSIZE4, RAMSIZE3, RAMSIZE2, RAMSIZE1, RAMSIZE0;
	input	BMSIZE3, BMSIZE2, BMSIZE1, BMSIZE0;
	input	WAIT2ND7, WAIT2ND6, WAIT2ND5, WAIT2ND4, WAIT2ND3, WAIT2ND2, WAIT2ND1, WAIT2ND0;
	input	PSELCPU, PSELBCD;
	input	CPUSTART/*, DECDYCUT*/;
	input	BASECKHS, RESB;
	input	SCANMODE;
	input	DFSIZE1, DFSIZE0;
	input	DFLEN;
	input	WED, FLSPM, GOFIRM;
	input	GATEAD1, GATEAD2, GATEAD3;
	input	CRCHLTEN;
// for EVA
        input   WAITFL2, ICEWAITMEM;
        input   SVI, SVVCOUT7, SVVCOUT6, SVVCOUT5, SVVCOUT4, SVVCOUT3, SVVCOUT2, SVVCOUT1, SVVCOUT0;
        input   ICECSGREGU, ICECSGREGA, ICEIFA4, ICEIFA3, ICEIFA2;
        input   ICEMSKNMI, ICEMSKDBG;
        // Ver1.51
        input   OCDMOD;
//
	wire	[19:0]	pc_inc;
// for EVA
//	wire	[7:0]	ID_stage1, ID_stage0, ID_stage1_dec;
	wire	[7:0]	ID_stage1_dec;
//
	wire	[7:0]	MEM_stage1, MEM_stage0;
// for EVA
//	wire	[1:0]	stage_adr;
//	wire	[14:0]	SP, sp_inc;
	wire	[14:0]	sp_inc;
//
	wire	[7:0]	A, X, B, C, D, E, H, L, buf1, buf0;
	wire	[7:0]	A_bank0,X_bank0,B_bank0,C_bank0,D_bank0,E_bank0,H_bank0,L_bank0;
	wire	[7:0]	A_bank1,X_bank1,B_bank1,C_bank1,D_bank1,E_bank1,H_bank1,L_bank1;
	wire	[7:0]	A_bank2,X_bank2,B_bank2,C_bank2,D_bank2,E_bank2,H_bank2,L_bank2;
	wire	[7:0]	A_bank3,X_bank3,B_bank3,C_bank3,D_bank3,E_bank3,H_bank3,L_bank3;
	wire	[3:0]	dec_alu_input10;
	wire	[3:0]	dec_alu_input20;
	wire	[3:0]	dec_alu_transout;
	wire	[4:0]	dec_alu_bitsh;
	wire	[3:0]	ES, CS, buf2;
// for EVA
//	wire	[15:0]	imdr;
//
	wire	[7:0]	PSW;
	wire	[1:0]	intisp;
	wire	[1:0]	BCDADJ;
	wire	[15:0]	ma_pre;
	wire		RVEON;

	wire		ivack, rstvec, skpack, dec_alu_add, dec_alu_sub, dec_alu_and, dec_alu_or, dec_alu_exor, dec_alu_ror;
	wire		dec_alu_rol, dec_alu_shr, dec_alu_shl, dec_alu_sar, dec_alu_mulu, dec_alu_carry, dec_word_access;
	wire		dec_alu_andbit, dec_alu_orbit, dec_alu_exorbit, dec_alu_biten; 
	wire		dec_xch_byte, dec_xchw_bc, dec_xchw_de, dec_xchw_hl, dec_SP_enable, dec_A_enable, dec_X_enable;
	wire		dec_B_enable, dec_C_enable, dec_D_enable, dec_E_enable, dec_H_enable, dec_L_enable, dec_ES_enable;
	wire		dec_Z_enable, dec_CY_enable, dec_AC_enable, dec_IE_enable, dec_ISP_enable, dec_NMIS_enable, dec_RBS_enable;
	wire		dec_buf0_enable, dec_buf1_enable, dec_buf2_enable, dec_ma_enable, dec_ma_data_sp, dec_ma_data_saddr_op1;
	wire		dec_ma_data_saddr_op2, dec_ma_data_sfr_op1, dec_ma_data_sfr_op2, dec_ma_data_op12, dec_ma_data_op23;
	wire		dec_ma_data_HL, dec_ma_data_HLop1, dec_ma_data_HLop2, dec_ma_data_HLB, dec_ma_data_HLC, dec_ma_data_DE;
	wire		dec_ma_data_DEop1, dec_ma_data_DEop2, dec_ma_data_SPop1, dec_ma_data_BCop12, dec_ma_data_Bop12, dec_ma_data_Cop12;
	wire		dec_sp_set_enable, dec_sp_inc, dec_sp_dec, dec_pc_inc1, dec_pc_inc2, dec_pc_inc3, dec_pc_inc4, dec_clear_stage;
	wire		dec_pc_set_enable, dec_pc_set_op01, dec_pc_set_op12, dec_pc_set_op123, dec_pc_set_AX, dec_pc_set_BC;
	wire		dec_pc_set_DE, dec_pc_set_HL, dec_pc_set_pc1, dec_pc_set_pc2, dec_pc_set_pc3, dec_pc_set_pc12, dec_pc_set_calt;
	wire		dec_pc_set_vec, dec_pc_set_brk, dec_pc_set_dbg, dec_pc_set_ret, dec_cpuwr_enable, dec_cpurd_enable;
	wire		dec_stage_cut_brtf, dec_stage_cut_ifbr, dec_ifbr_not, dec_ifbr_zero, dec_ifbr_ht;
	wire		dec_mem_stage_op2, dec_mem_stage_op3, dec_mem_stage_op23, dec_set_buf_retadr, dec_set_buf_intr;
	wire		dec_skc, dec_sknc, dec_skz, dec_sknz, dec_skh, dec_sknh, dec_prefix, dec_halt, dec_stop;
	wire		dec_movs, dec_cmps, CPUEN, slreg, slmirr, maw1, stage_cut, MAA, A_access, X_access, B_access, C_access;
	wire		D_access, E_access, H_access, L_access, INT_access, skp_block, intblock, PSW_block, SP_enable, CS_enable;
	wire		stage_cut_br, pc_set_brk, pc_set_dbg, waitdma, ivack_pre, fchiram, fchiram_skp, romrd_skp;
	wire		pc_wait_flg, stby_wait_flg, reg_wait, pa_data_buf, pa_data_mem, pa_data_spen, pa_st2;
	wire		data_hazard_flg, data_hazard, sp_hazard, pswlock;
	wire		wait_block_brtf, pswen, INT_wait, dopen, waitint, prefix_ack;
	wire		exmmsk, flmask, mem_access, stbst;
	wire		dec_alu_transin, cpuwr_reg, wait2ndsfr, sl2ndwait_pre;
// for EVA
	wire	[14:0]	SP_usr, SP_sv;
	wire		dec_alt1, dec_alt2, svmodi;
//
	wire	[3:0]	dec_alu_input10_dmy;
	wire		waitdflash, sldfwait_pre;
	wire		GATEAD1, GATEAD2, GATEAD3;
	wire		CRCHLTEN;

	assign dec_alu_input10_dmy[3] = dec_alu_input10[3];
	assign dec_alu_input10_dmy[2] = dec_alu_input10[2] ^ (dec_alu_input10[3] & ~dec_alu_input10[2] & dec_alu_input10[1] & dec_alu_input10[0]) ;
	assign dec_alu_input10_dmy[1] = dec_alu_input10[1];
	assign dec_alu_input10_dmy[0] = dec_alu_input10[0] ^ (dec_alu_input10[3] & ~dec_alu_input10[2] & dec_alu_input10[1] & dec_alu_input10[0]) ;

	QLK0RCPUEVA0V3_DEC dec(
// for EVA
//		.ID_stage1(ID_stage1_dec), .ID_stage0(ID_stage0), .decout_mask_reg(decout_mask_reg),
		.ID_stage1(ID_stage1_dec), 
                .ID_stage0({IDADR7, IDADR6, IDADR5, IDADR4, IDADR3, IDADR2, IDADR1, IDADR0}),
//
// for EVA
//		.stage_adr(stage_adr), .ivack(ivack),  .rstvec(rstvec), .skpack(skpack),
                .stage_adr({STAGEADR1, STAGEADR0}), .ivack(ivack), .rstvec(rstvec), .skpack(skpack),
//
		.dec_alu_input10(dec_alu_input10), .dec_alu_input20(dec_alu_input20),
		.dec_alu_add(dec_alu_add), .dec_alu_sub(dec_alu_sub), .dec_alu_and(dec_alu_and),
		.dec_alu_or(dec_alu_or), .dec_alu_exor(dec_alu_exor),
		.dec_alu_andbit(dec_alu_andbit), .dec_alu_orbit(dec_alu_orbit), .dec_alu_exorbit(dec_alu_exorbit),
		.dec_alu_ror(dec_alu_ror), .dec_alu_rol(dec_alu_rol),
		.dec_alu_shr(dec_alu_shr), .dec_alu_shl(dec_alu_shl), .dec_alu_sar(dec_alu_sar),
		.dec_alu_mulu(dec_alu_mulu), .dec_alu_carry(dec_alu_carry),
		.dec_alu_transin(dec_alu_transin), .dec_alu_transout(dec_alu_transout),
		.dec_alu_bitsh(dec_alu_bitsh), .dec_alu_biten(dec_alu_biten),
		.dec_word_access(dec_word_access),
		.dec_xch_byte(dec_xch_byte), .dec_xchw_bc(dec_xchw_bc), 
		.dec_xchw_de(dec_xchw_de), .dec_xchw_hl(dec_xchw_hl), 
		.dec_SP_enable(dec_SP_enable),
		.dec_A_enable(dec_A_enable), .dec_X_enable(dec_X_enable),
		.dec_B_enable(dec_B_enable), .dec_C_enable(dec_C_enable),
		.dec_D_enable(dec_D_enable), .dec_E_enable(dec_E_enable),
		.dec_H_enable(dec_H_enable), .dec_L_enable(dec_L_enable),
		.dec_ES_enable(dec_ES_enable),
		.dec_Z_enable(dec_Z_enable), .dec_CY_enable(dec_CY_enable),
		.dec_AC_enable(dec_AC_enable), .dec_IE_enable(dec_IE_enable),
		.dec_ISP_enable(dec_ISP_enable), .dec_NMIS_enable(dec_NMIS_enable), .dec_RBS_enable(dec_RBS_enable),
		.dec_buf0_enable(dec_buf0_enable), .dec_buf1_enable(dec_buf1_enable), .dec_buf2_enable(dec_buf2_enable),
		.dec_ma_enable(dec_ma_enable),
		.dec_ma_data_sp(dec_ma_data_sp),
		.dec_ma_data_saddr_op1(dec_ma_data_saddr_op1), .dec_ma_data_saddr_op2(dec_ma_data_saddr_op2),
		.dec_ma_data_sfr_op1(dec_ma_data_sfr_op1), .dec_ma_data_sfr_op2(dec_ma_data_sfr_op2),
		.dec_ma_data_op12(dec_ma_data_op12), .dec_ma_data_op23(dec_ma_data_op23),
		.dec_ma_data_HL(dec_ma_data_HL), .dec_ma_data_HLop1(dec_ma_data_HLop1), .dec_ma_data_HLop2(dec_ma_data_HLop2),
		.dec_ma_data_HLB(dec_ma_data_HLB), .dec_ma_data_HLC(dec_ma_data_HLC),
		.dec_ma_data_DE(dec_ma_data_DE), .dec_ma_data_DEop1(dec_ma_data_DEop1), .dec_ma_data_DEop2(dec_ma_data_DEop2),
		.dec_ma_data_SPop1(dec_ma_data_SPop1),
		.dec_ma_data_BCop12(dec_ma_data_BCop12),
		.dec_ma_data_Bop12(dec_ma_data_Bop12), .dec_ma_data_Cop12(dec_ma_data_Cop12),
		.dec_sp_set_enable(dec_sp_set_enable), .dec_sp_inc(dec_sp_inc), .dec_sp_dec(dec_sp_dec),
		.dec_pc_inc1(dec_pc_inc1), .dec_pc_inc2(dec_pc_inc2),
		.dec_pc_inc3(dec_pc_inc3), .dec_pc_inc4(dec_pc_inc4),
		.dec_clear_stage(dec_clear_stage), .dec_pc_set_enable(dec_pc_set_enable),
		.dec_pc_set_op01(dec_pc_set_op01), .dec_pc_set_op12(dec_pc_set_op12), .dec_pc_set_op123(dec_pc_set_op123),
		.dec_pc_set_AX(dec_pc_set_AX), .dec_pc_set_BC(dec_pc_set_BC),
		.dec_pc_set_DE(dec_pc_set_DE), .dec_pc_set_HL(dec_pc_set_HL),
		.dec_pc_set_pc1(dec_pc_set_pc1), .dec_pc_set_pc2(dec_pc_set_pc2), .dec_pc_set_pc3(dec_pc_set_pc3),
		.dec_pc_set_pc12(dec_pc_set_pc12),
		.dec_pc_set_calt(dec_pc_set_calt), .dec_pc_set_vec(dec_pc_set_vec),
		.dec_pc_set_brk(dec_pc_set_brk), .dec_pc_set_dbg(dec_pc_set_dbg),
		.dec_pc_set_ret(dec_pc_set_ret),
		.dec_cpuwr_enable(dec_cpuwr_enable), .dec_cpurd_enable(dec_cpurd_enable),
		.dec_stage_cut_brtf(dec_stage_cut_brtf), .dec_stage_cut_ifbr(dec_stage_cut_ifbr),
		.dec_ifbr_not(dec_ifbr_not), .dec_ifbr_zero(dec_ifbr_zero), .dec_ifbr_ht(dec_ifbr_ht),
		.dec_mem_stage_op2(dec_mem_stage_op2), .dec_mem_stage_op3(dec_mem_stage_op3), .dec_mem_stage_op23(dec_mem_stage_op23),
		.dec_set_buf_retadr(dec_set_buf_retadr), .dec_set_buf_intr(dec_set_buf_intr),
		.dec_skc(dec_skc), .dec_sknc(dec_sknc), .dec_skz(dec_skz), .dec_sknz(dec_sknz), .dec_skh(dec_skh), .dec_sknh(dec_sknh),
		.dec_prefix(dec_prefix), .dec_halt(dec_halt), .dec_stop(dec_stop), .dec_movs(dec_movs), .dec_cmps(dec_cmps),
// for EVA
		.dec_alt1(dec_alt1), .dec_alt2(dec_alt2),
//
		.cpuen(CPUEN), .baseck(BASECKHS), .resb(RESB), .scanmode(SCANMODE) );

	QLK0RCPUEVA0V3_ALU alu(
// for EVA
//		.imdr(imdr), .pselcpu(PSELCPU),  .pselbcd(PSELBCD), .slreg(slreg), .slmirr(slmirr),
                .pselcpu(PSELCPU),  .pselbcd(PSELBCD), .slreg(slreg), .slmirr(slmirr),
                .imdr({IMDR15, IMDR14, IMDR13, IMDR12, IMDR11, IMDR10, IMDR9, IMDR8,
                       IMDR7, IMDR6, IMDR5, IMDR4, IMDR3, IMDR2, IMDR1, IMDR0}),
//
		.vpa({MA3, MA2, MA1, MA0}),
		.pid({PID31, PID30, PID29, PID28, PID27, PID26, PID25, PID24, PID23, PID22, PID21, PID20, PID19, PID18, PID17, PID16,
		      PID15, PID14, PID13, PID12, PID11, PID10, PID9, PID8, PID7, PID6, PID5, PID4, PID3, PID2, PID1, PID0}),
		.mdw({MDW15, MDW14, MDW13, MDW12, MDW11, MDW10, MDW9, MDW8, MDW7, MDW6, MDW5, MDW4, MDW3, MDW2, MDW1, MDW0}),
		.biten({BITEN7, BITEN6, BITEN5, BITEN4, BITEN3, BITEN2, BITEN1, BITEN0}),
		.pc({PC19, PC18, PC17, PC16, PC15, PC14, PC13, PC12, PC11, PC10, PC9, PC8, PC7, PC6, PC5, PC4, PC3, PC2, PC1, PC0}),
		.ma_pre(ma_pre), .maw1(maw1), .pc_inc(pc_inc), .wdop(WDOP), .wdwr(WDWR),
// for EVA
//		.ID_stage0(ID_stage0), .MEM_stage0(MEM_stage0), .MEM_stage1(MEM_stage1),
		.ID_stage0({IDADR7, IDADR6, IDADR5, IDADR4, IDADR3, IDADR2, IDADR1, IDADR0}),
		.MEM_stage0(MEM_stage0), .MEM_stage1(MEM_stage1),
//
		.cpuwr(CPUWR), .cpuwr_reg(cpuwr_reg), .cpurd(CPURD), .stage_cut(stage_cut),
		.A(A), .X(X), .B(B), .C(C), .D(D), .E(E), .H(H), .L(L), .CS(CS), .ES(ES), .PSW(PSW), .MAA(MAA), .BCDADJ(BCDADJ),
		.A_bank0(A_bank0), .X_bank0(X_bank0), .B_bank0(B_bank0), .C_bank0(C_bank0),
		.D_bank0(D_bank0), .E_bank0(E_bank0), .H_bank0(H_bank0), .L_bank0(L_bank0),
		.A_bank1(A_bank1), .X_bank1(X_bank1), .B_bank1(B_bank1), .C_bank1(C_bank1),
		.D_bank1(D_bank1), .E_bank1(E_bank1), .H_bank1(H_bank1), .L_bank1(L_bank1),
		.A_bank2(A_bank2), .X_bank2(X_bank2), .B_bank2(B_bank2), .C_bank2(C_bank2),
		.D_bank2(D_bank2), .E_bank2(E_bank2), .H_bank2(H_bank2), .L_bank2(L_bank2),
		.A_bank3(A_bank3), .X_bank3(X_bank3), .B_bank3(B_bank3), .C_bank3(C_bank3),
		.D_bank3(D_bank3), .E_bank3(E_bank3), .H_bank3(H_bank3), .L_bank3(L_bank3),
		.A_access(A_access), .X_access(X_access), .B_access(B_access), .C_access(C_access),
		.D_access(D_access), .E_access(E_access), .H_access(H_access), .L_access(L_access),
		.INT_access(INT_access), .skp_block(skp_block),
		.intblock(intblock), .PSW_block(PSW_block), .SP_enable(SP_enable), .CS_enable(CS_enable),
		.stage_cut_br(stage_cut_br), .pc_set_brk(pc_set_brk), .pc_set_dbg(pc_set_dbg),
// for EVA
//		.buf2(buf2), .buf1(buf1), .buf0(buf0), .SP(SP), .sp_inc(sp_inc),
		.buf2(buf2), .buf1(buf1), .buf0(buf0), .sp_inc(sp_inc),
                .SP({SP15, SP14, SP13, SP12, SP11, SP10, SP9, SP8, SP7, SP6, SP5, SP4, SP3, SP2, SP1}), .SP0(SP0),
//
		.dmard(DMARD), .dmawr(DMAWR), .dmawdop(DMAWDOP), .waitdma(waitdma),
		.ivack(ivack), .ivack_pre(ivack_pre), .intisp(intisp),
		.fchiram(fchiram), .fchiram_skp(fchiram_skp), .romrd_skp(romrd_skp),
		.pc_wait_flg(pc_wait_flg), .reg_wait(reg_wait),
		.pa_data_buf(pa_data_buf), .pa_data_mem(pa_data_mem), .pa_data_spen(pa_data_spen),
		.pa_st2(pa_st2), .slflash(SLFLASH),
		.data_hazard_flg(data_hazard_flg), .data_hazard(data_hazard), .sp_hazard(sp_hazard),
		.dec_alu_input10(dec_alu_input10_dmy), .dec_alu_input20(dec_alu_input20),
		.dec_alu_add(dec_alu_add), .dec_alu_sub(dec_alu_sub), .dec_alu_and(dec_alu_and),
		.dec_alu_or(dec_alu_or), .dec_alu_exor(dec_alu_exor),
		.dec_alu_andbit(dec_alu_andbit), .dec_alu_orbit(dec_alu_orbit), .dec_alu_exorbit(dec_alu_exorbit),
		.dec_alu_ror(dec_alu_ror), .dec_alu_rol(dec_alu_rol),
		.dec_alu_shr(dec_alu_shr), .dec_alu_shl(dec_alu_shl), .dec_alu_sar(dec_alu_sar),
		.dec_alu_mulu(dec_alu_mulu), .dec_alu_carry(dec_alu_carry),
		.dec_alu_transin(dec_alu_transin), .dec_alu_transout(dec_alu_transout),
		.dec_alu_bitsh(dec_alu_bitsh), .dec_alu_biten(dec_alu_biten),
		.dec_word_access(dec_word_access),
		.dec_xch_byte(dec_xch_byte), .dec_xchw_bc(dec_xchw_bc),
		.dec_xchw_de(dec_xchw_de), .dec_xchw_hl(dec_xchw_hl),
		.dec_A_enable(dec_A_enable), .dec_X_enable(dec_X_enable),
		.dec_B_enable(dec_B_enable), .dec_C_enable(dec_C_enable),
		.dec_D_enable(dec_D_enable), .dec_E_enable(dec_E_enable),
		.dec_H_enable(dec_H_enable), .dec_L_enable(dec_L_enable),
		.dec_ES_enable(dec_ES_enable),
		.dec_Z_enable(dec_Z_enable), .dec_CY_enable(dec_CY_enable),
		.dec_AC_enable(dec_AC_enable), .dec_IE_enable(dec_IE_enable),
		.dec_ISP_enable(dec_ISP_enable), .dec_RBS_enable(dec_RBS_enable),
		.dec_buf0_enable(dec_buf0_enable), .dec_buf1_enable(dec_buf1_enable), .dec_buf2_enable(dec_buf2_enable),
		.dec_SP_enable(dec_SP_enable),
		.dec_cpuwr_enable(dec_cpuwr_enable),
		.dec_cpurd_enable(dec_cpurd_enable),
		.dec_sp_set_enable(dec_sp_set_enable), .dec_sp_inc(dec_sp_inc),  .dec_sp_dec(dec_sp_dec),
		.dec_stage_cut_brtf(dec_stage_cut_brtf), .dec_stage_cut_ifbr(dec_stage_cut_ifbr),
		.dec_ifbr_not(dec_ifbr_not), .dec_ifbr_zero(dec_ifbr_zero), .dec_ifbr_ht(dec_ifbr_ht),
		.dec_set_buf_retadr(dec_set_buf_retadr), .dec_set_buf_intr(dec_set_buf_intr),
		.dec_skc(dec_skc), .dec_sknc(dec_sknc), .dec_skz(dec_skz), .dec_sknz(dec_sknz),
		.dec_skh(dec_skh), .dec_sknh(dec_sknh),
		.dec_movs(dec_movs), .dec_cmps(dec_cmps),
		.dec_ma_enable(dec_ma_enable),
		.skpack(skpack), .skipexe(SKIPEXE), .pswlock(pswlock),
		.wait_block_brtf(wait_block_brtf),
		.mem_access(mem_access),
// for EVA
                .SP_usr(SP_usr), .SP_sv(SP_sv),
                .svmod(SVMOD), .svmodi(svmodi),
                .alt1(ALT1), .alt2(ALT2),
                .spinc(SPINC), .spdec(SPDEC),
                .icecsgregu(ICECSGREGU), .icecsgrega(ICECSGREGA), .iceifa({ICEIFA4, ICEIFA3, ICEIFA2}),
                .icedo({ICEDO31, ICEDO30, ICEDO29, ICEDO28, ICEDO27, ICEDO26, ICEDO25, ICEDO24,ICEDO23,
                        ICEDO22, ICEDO21, ICEDO20, ICEDO19, ICEDO18, ICEDO17, ICEDO16,ICEDO15,
                        ICEDO14, ICEDO13, ICEDO12, ICEDO11, ICEDO10, ICEDO9, ICEDO8,
                        ICEDO7, ICEDO6, ICEDO5, ICEDO4, ICEDO3, ICEDO2, ICEDO1, ICEDO0}),
//
		.cpuen(CPUEN), .pswen(pswen), .baseck(BASECKHS), .resb(RESB), .scanmode(SCANMODE),
		.RVEON(RVEON)
		);

	QLK0RCPUEVA0V3_ADR adr(
// for EVA
//		.ID_stage1(ID_stage1), .ID_stage0(ID_stage0), .ID_stage1_dec(ID_stage1_dec),
                .ID_stage1_dec(ID_stage1_dec),
                .ID_stage3({IDADR31, IDADR30, IDADR29, IDADR28, IDADR27, IDADR26, IDADR25, IDADR24}),
                .ID_stage2({IDADR23, IDADR22, IDADR21, IDADR20, IDADR19, IDADR18, IDADR17, IDADR16}),
                .ID_stage1({IDADR15, IDADR14, IDADR13, IDADR12, IDADR11, IDADR10, IDADR9, IDADR8}),
                .ID_stage0({IDADR7, IDADR6, IDADR5, IDADR4, IDADR3, IDADR2, IDADR1, IDADR0}),
//
		.MEM_stage1(MEM_stage1), .MEM_stage0(MEM_stage0),
// for EVA
//		.stage_adr(stage_adr), .pc_inc(pc_inc),
                .stage_adr({STAGEADR1, STAGEADR0}), .pc_inc(pc_inc),
//
		.pc_wait_flg(pc_wait_flg), .stby_wait_flg(stby_wait_flg), .reg_wait(reg_wait),
		.pa_data_buf(pa_data_buf), .pa_data_mem(pa_data_mem), .pa_st2(pa_st2), .pa_data_spen(pa_data_spen),
		.pa({PA19, PA18, PA17, PA16, PA15, PA14, PA13, PA12, PA11, PA10, PA9, PA8, PA7, PA6, PA5, PA4, PA3, PA2}),
		.pc({PC19, PC18, PC17, PC16, PC15, PC14, PC13, PC12, PC11, PC10, PC9, PC8, PC7, PC6, PC5, PC4, PC3, PC2, PC1, PC0}),
		.pid({PID31, PID30, PID29, PID28, PID27, PID26, PID25, PID24, PID23, PID22, PID21, PID20, PID19, PID18, PID17, PID16,
		      PID15, PID14, PID13, PID12, PID11, PID10, PID9, PID8, PID7, PID6, PID5, PID4, PID3, PID2, PID1, PID0}),
		.data_hazard_flg(data_hazard_flg), .data_hazard(data_hazard), .sp_hazard(sp_hazard),
		.A_access(A_access), .X_access(X_access), .B_access(B_access), .C_access(C_access),
		.D_access(D_access), .E_access(E_access), .H_access(H_access), .L_access(L_access),
		.dec_RBS_enable(dec_RBS_enable),
		.INT_access(INT_access), .INT_wait(INT_wait), .wait2ndsfr(wait2ndsfr), .sl2ndwait_pre(sl2ndwait_pre), .dopen(dopen),
		.dec_NMIS_enable(dec_NMIS_enable), .SP_enable(SP_enable),
		.CS_enable(CS_enable),
		.dec_SP_enable(dec_SP_enable),
		.dec_pc_inc1(dec_pc_inc1), .dec_pc_inc2(dec_pc_inc2),
		.dec_pc_inc3(dec_pc_inc3), .dec_pc_inc4(dec_pc_inc4),
		.dec_clear_stage(dec_clear_stage), .dec_pc_set_enable(dec_pc_set_enable),
		.dec_pc_set_op01(dec_pc_set_op01), .dec_pc_set_op12(dec_pc_set_op12), .dec_pc_set_op123(dec_pc_set_op123),
		.dec_pc_set_AX(dec_pc_set_AX), .dec_pc_set_BC(dec_pc_set_BC),
		.dec_pc_set_DE(dec_pc_set_DE), .dec_pc_set_HL(dec_pc_set_HL),
		.dec_pc_set_pc1(dec_pc_set_pc1), .dec_pc_set_pc2(dec_pc_set_pc2), .dec_pc_set_pc3(dec_pc_set_pc3),
		.dec_pc_set_pc12(dec_pc_set_pc12),
		.dec_pc_set_calt(dec_pc_set_calt), .dec_pc_set_vec(dec_pc_set_vec),
		.dec_pc_set_brk(dec_pc_set_brk), .dec_pc_set_dbg(dec_pc_set_dbg),
		.dec_pc_set_ret(dec_pc_set_ret),
		.dec_ma_enable(dec_ma_enable),
		.dec_ma_data_sp(dec_ma_data_sp),
		.dec_ma_data_saddr_op1(dec_ma_data_saddr_op1), .dec_ma_data_saddr_op2(dec_ma_data_saddr_op2),
		.dec_ma_data_sfr_op1(dec_ma_data_sfr_op1), .dec_ma_data_sfr_op2(dec_ma_data_sfr_op2),
		.dec_ma_data_op12(dec_ma_data_op12), .dec_ma_data_op23(dec_ma_data_op23),
		.dec_ma_data_HL(dec_ma_data_HL), .dec_ma_data_HLop1(dec_ma_data_HLop1), .dec_ma_data_HLop2(dec_ma_data_HLop2),
		.dec_ma_data_HLB(dec_ma_data_HLB), .dec_ma_data_HLC(dec_ma_data_HLC),
		.dec_ma_data_DE(dec_ma_data_DE), .dec_ma_data_DEop1(dec_ma_data_DEop1), .dec_ma_data_DEop2(dec_ma_data_DEop2),
		.dec_ma_data_SPop1(dec_ma_data_SPop1),
		.dec_ma_data_BCop12(dec_ma_data_BCop12),
		.dec_ma_data_Bop12(dec_ma_data_Bop12), .dec_ma_data_Cop12(dec_ma_data_Cop12),
		.dec_sp_set_enable(dec_sp_set_enable), .dec_cpurd_enable(dec_cpurd_enable), .dec_cpuwr_enable(dec_cpuwr_enable),
		.dec_mem_stage_op2(dec_mem_stage_op2), .dec_mem_stage_op3(dec_mem_stage_op3), .dec_mem_stage_op23(dec_mem_stage_op23),
		.dec_prefix(dec_prefix), .stage_cut(stage_cut),
		.A(A), .X(X), .B(B), .C(C), .D(D), .E(E), .H(H), .L(L), .CS(CS), .ES(ES),
		.buf2(buf2), .buf1(buf1), .buf0(buf0),
		.ma({MA15, MA14, MA13, MA12, MA11, MA10, MA9, MA8, MA7, MA6, MA5, MA4, MA3, MA2, MA1, MA0}),
		.ma_pre(ma_pre), .maw1(maw1),
		.exma({EXMA3, EXMA2, EXMA1, EXMA0}),
		.slmem(SLMEM), .slflash(SLFLASH), .slreg(slreg), .slmirr(slmirr), .slexm(SLEXM), .slbmem(SLBMEM), .sliram(SLIRAM),
		.cpuwr(CPUWR), .cpuwr_reg(cpuwr_reg), .cpurd(CPURD),
// for EVA
//		.imdr(imdr),
                .imdr({IMDR15, IMDR14, IMDR13, IMDR12, IMDR11, IMDR10, IMDR9, IMDR8,
                       IMDR7, IMDR6, IMDR5, IMDR4, IMDR3, IMDR2, IMDR1, IMDR0}),
//
		.dmama({DMAMA15, DMAMA14, DMAMA13, DMAMA12, DMAMA11, DMAMA10, DMAMA9, DMAMA8, DMAMA7, DMAMA6, DMAMA5,
			DMAMA4, DMAMA3, DMAMA2, DMAMA1, DMAMA0}),
		.hltst(HLTST), .stbst(stbst), .dmarq(DMARQ), .dmaack(DMAACK), .waitdma(waitdma), .waitint(waitint),
		.waitfl(WAITFL), .waitexm(WAITEXM), .waitmod(WAITMOD), .waitmem(WAITMEM),
		.vcout({VCOUT6, VCOUT5, VCOUT4, VCOUT3, VCOUT2, VCOUT1}),
// for EVA
//		.MAA(MAA), .IE(PSW[7]), .SP(SP), .sp_inc(sp_inc), .wdop(WDOP),
                .MAA(MAA), .IE(PSW[7]), .sp_inc(sp_inc), .wdop(WDOP),
                .SP({SP15, SP14, SP13, SP12, SP11, SP10, SP9, SP8, SP7, SP6, SP5, SP4, SP3, SP2, SP1}),
//
		.intdbg(INTDBG), .intnmi(INTNMI), .intrq3(INTRQ3), .intrq2(INTRQ2), .intrq1(INTRQ1), .intrq0(INTRQ0),
		.isp(PSW[2:1]), .intack(INTACK), .ivack(ivack), .ivack_pre(ivack_pre), .monmd(MONMD), .monmdstp(MONMDSTP), .softbrk(SOFTBRK),
		.intisp(intisp), .intblock(intblock), .PSW_block(PSW_block), .skp_block(skp_block),  .wait_block_brtf(wait_block_brtf),
		.stage_cut_br(stage_cut_br), .pc_set_brk(pc_set_brk), .pc_set_dbg(pc_set_dbg),
		.prefix_ack(prefix_ack), .fchiram(fchiram), .fchiram_skp(fchiram_skp), .romrd_skp(romrd_skp), .rstvec(rstvec),
		.flsize({FLSIZE3, FLSIZE2, FLSIZE1, FLSIZE0}), .bfsize({BFSIZE3, BFSIZE2, BFSIZE1, BFSIZE0}),
		.ramsize({RAMSIZE7, RAMSIZE6, RAMSIZE5, RAMSIZE4, RAMSIZE3, RAMSIZE2, RAMSIZE1, RAMSIZE0}),
		.bmsize({BMSIZE3, BMSIZE2, BMSIZE1, BMSIZE0}),
		.wait2nd({WAIT2ND7, WAIT2ND6, WAIT2ND5, WAIT2ND4, WAIT2ND3, WAIT2ND2, WAIT2ND1, WAIT2ND0}),
		.exmmsk(exmmsk), .flmask(flmask), /*.decdycut(DECDYCUT),*/ .brkmsk(BRKMSK),
		.flread(FLREAD), .fchram(FCHRAM), .mem_access(mem_access),
// for EVA
                .svi(SVI), .svvcout({SVVCOUT7, SVVCOUT6, SVVCOUT5, SVVCOUT4, SVVCOUT3, SVVCOUT2, SVVCOUT1, SVVCOUT0}),
                .svintack(SVINTACK), .svmod(SVMOD), .svmodf(SVMODF), .svmodi(svmodi),
                .dec_alt1(dec_alt1), .dec_alt2(dec_alt2), .alt1(ALT1), .alt2(ALT2),
                .dec_sp_inc(dec_sp_inc), .idpop(IDPOP),
                .flreadb({FLREADB3, FLREADB2, FLREADB1, FLREADB0}),
                .prefix(PREFIX), .pcwaitf(PCWAITF),
                .icemsknmi(ICEMSKNMI), .icemskdbg(ICEMSKDBG),
                .cpumisal(CPUMISAL), .sprel(SPREL),
                .pswen(pswen),
                // Ver1.51
                .ocdmod(OCDMOD),
//
		.cpuen(CPUEN), .baseck(BASECKHS), .resb(RESB), .scanmode(SCANMODE),
		.dfsize({DFSIZE1,DFSIZE0}), .dflen(DFLEN),
		.sldflash(SLDFLASH), .drdclk(DRDCLK), .waitdflash(waitdflash), .sldfwait_pre(sldfwait_pre),
		.wed(WED), .flspm(FLSPM), .gofirm(GOFIRM),
		.RVEON(RVEON), 
		.gatead1(GATEAD1), .gatead2(GATEAD2), .gatead3(GATEAD3),
		.mdw({MDW15, MDW14, MDW13, MDW12, MDW11, MDW10, MDW9, MDW8, MDW7, MDW6, MDW5, MDW4, MDW3, MDW2, MDW1, MDW0}),
		.monpc({MONPC19, MONPC18, MONPC17, MONPC16, MONPC15, MONPC14, MONPC13, MONPC12, MONPC11, MONPC10, 
			MONPC9, MONPC8, MONPC7, MONPC6, MONPC5, MONPC4, MONPC3, MONPC2, MONPC1, MONPC0}),
		.monma({MONMA15, MONMA14, MONMA13, MONMA12, MONMA11, MONMA10, 
			MONMA9, MONMA8, MONMA7, MONMA6, MONMA5, MONMA4, MONMA3, MONMA2, MONMA1, MONMA0}),
		.monmdr({MONMDR15, MONMDR14, MONMDR13, MONMDR12, MONMDR11, MONMDR10, 
			 MONMDR9, MONMDR8, MONMDR7, MONMDR6, MONMDR5, MONMDR4, MONMDR3, MONMDR2, MONMDR1, MONMDR0}),
		.monmdw({MONMDW15, MONMDW14, MONMDW13, MONMDW12, MONMDW11, MONMDW10, 
			 MONMDW9, MONMDW8, MONMDW7, MONMDW6, MONMDW5, MONMDW4, MONMDW3, MONMDW2, MONMDW1, MONMDW0})
		);

	QLK0RCPUEVA0V3_CLK clk(
		.mdr({MDR15, MDR14, MDR13, MDR12, MDR11, MDR10, MDR9, MDR8, MDR7, MDR6, MDR5, MDR4, MDR3, MDR2, MDR1, MDR0}),
// for EVA
//		.imdr(imdr), .pselcpu(PSELCPU), .pselbcd(PSELBCD), .slreg(slreg), .rga(MA4), .vpa({MA3, MA2, MA1, MA0}),
                .pselcpu(PSELCPU), .pselbcd(PSELBCD), .slreg(slreg), .rga(MA4), .vpa({MA3, MA2, MA1, MA0}),
                .imdr({IMDR15, IMDR14, IMDR13, IMDR12, IMDR11, IMDR10, IMDR9, IMDR8,
                       IMDR7, IMDR6, IMDR5, IMDR4, IMDR3, IMDR2, IMDR1, IMDR0}),
//
		.dec_set_buf_retadr(dec_set_buf_retadr), .dec_set_buf_intr(dec_set_buf_intr),
		.dec_halt(dec_halt), .dec_stop(dec_stop), .stben(STBEN), .pc_wait_flg(pc_wait_flg),
		.stby_wait_flg(stby_wait_flg),
		.intdbg(INTDBG), .intnmi(INTNMI), .intrq3(INTRQ3), .intrq2(INTRQ2), .intrq1(INTRQ1), .intrq0(INTRQ0),
		.cpurd(CPURD), .wdop(WDOP),
// for EVA
//		.SP(SP), .PSW(PSW), .CS(CS), .ES(ES), .MAA(MAA), .BCDADJ(BCDADJ),
                .PSW(PSW), .CS(CS), .ES(ES), .MAA(MAA), .BCDADJ(BCDADJ),
                .SP({SP15, SP14, SP13, SP12, SP11, SP10, SP9, SP8, SP7, SP6, SP5, SP4, SP3, SP2, SP1}),
//
		.A_bank0(A_bank0), .X_bank0(X_bank0), .B_bank0(B_bank0), .C_bank0(C_bank0),
		.D_bank0(D_bank0), .E_bank0(E_bank0), .H_bank0(H_bank0), .L_bank0(L_bank0),
		.A_bank1(A_bank1), .X_bank1(X_bank1), .B_bank1(B_bank1), .C_bank1(C_bank1),
		.D_bank1(D_bank1), .E_bank1(E_bank1), .H_bank1(H_bank1), .L_bank1(L_bank1),
		.A_bank2(A_bank2), .X_bank2(X_bank2), .B_bank2(B_bank2), .C_bank2(C_bank2),
		.D_bank2(D_bank2), .E_bank2(E_bank2), .H_bank2(H_bank2), .L_bank2(L_bank2),
		.A_bank3(A_bank3), .X_bank3(X_bank3), .B_bank3(B_bank3), .C_bank3(C_bank3),
		.D_bank3(D_bank3), .E_bank3(E_bank3), .H_bank3(H_bank3), .L_bank3(L_bank3),
		.INT_wait(INT_wait), .wait2ndsfr(wait2ndsfr), .sl2ndwait_pre(sl2ndwait_pre), .waitdma(waitdma), .waitint(waitint),
		.dmarq(DMARQ), .dopen(dopen), .dmaack(DMAACK),
		.waitfl(WAITFL), .waitmod(WAITMOD), .waitexm(WAITEXM), .dmaen(DMAEN), .dmawait(DMAWAIT), .ocdwait(OCDWAIT),
		.pswlock(pswlock), .exmmsk(exmmsk), .flmask(flmask), .hltst(HLTST), .stpst(STPST), .stbst(stbst),
// for EVA
                .SP_usr(SP_usr), .SP_sv(SP_sv), .svmod(SVMOD), .alt1(ALT1),
                .svi(SVI),
                .waitfl2(WAITFL2), .icewaitmem(ICEWAITMEM),
                .cpumask(CPUMASK),
//
		.cpustart(CPUSTART), .cpuen(CPUEN), .pswen(pswen), .baseck(BASECKHS), .resb(RESB), .scanmode(SCANMODE),
		.sldfwait_pre(sldfwait_pre), .waitdflash(waitdflash),
		.RVEON(RVEON), .crchlten(CRCHLTEN)
		);

endmodule

/********************************************************************************/
/* K0R EVA ADR Block                                                           	*/
/*                                                          Made K.Tanaka       */
/********************************************************************************/
/* Ver1.00  New                                                                 */
/* Ver1.50  Add flread                                2007.05.30 K.Tanaka       */
/*              fchram                                2007.05.30 K.Tanaka       */
/*              mem_access                            2007.05.30 K.Tanaka       */
/*              stbst                                 2007.07.02 K.Tanaka       */
/* Ver1.51  Add ocdmod                                2007.11.30 K.Tanaka       */
/* Ver1.52  Modified MONMD Signal during svmod        2008.02.26 K.Tanaka       */
/* Ver2.01  Modified CPUMISAL Signal                  2008.08.29 K.Tanaka       */
/********************************************************************************/
module QLK0RCPUEVA0V3_ADR(
	ID_stage1, ID_stage0, ID_stage1_dec, 
	MEM_stage1, MEM_stage0,
	stage_adr, pc, pc_inc, pc_wait_flg, stby_wait_flg, reg_wait,
	pa_data_buf, pa_data_mem, pa_data_spen,
	pa_st2, pa, pid, data_hazard_flg, data_hazard, sp_hazard,
	dec_NMIS_enable, SP_enable,
	CS_enable,
	A_access, X_access, B_access, C_access,
	D_access, E_access, H_access, L_access,
	dec_RBS_enable, INT_access, INT_wait, wait2ndsfr, sl2ndwait_pre, dopen,
	dec_SP_enable,
	dec_pc_inc1, dec_pc_inc2, dec_pc_inc3, dec_pc_inc4,
	dec_clear_stage, dec_pc_set_enable,
	dec_pc_set_op01, dec_pc_set_op12, dec_pc_set_op123,
	dec_pc_set_AX, dec_pc_set_BC,
	dec_pc_set_DE, dec_pc_set_HL,
	dec_pc_set_pc1, dec_pc_set_pc2, dec_pc_set_pc3,
	dec_pc_set_pc12,
	dec_pc_set_calt, dec_pc_set_vec,
	dec_pc_set_brk, dec_pc_set_dbg,
	dec_pc_set_ret,
	dec_ma_enable,
	dec_ma_data_sp,
	dec_ma_data_saddr_op1, dec_ma_data_saddr_op2,
	dec_ma_data_sfr_op1, dec_ma_data_sfr_op2,
	dec_ma_data_op12, dec_ma_data_op23,
	dec_ma_data_HL, dec_ma_data_HLop1, dec_ma_data_HLop2,
	dec_ma_data_HLB, dec_ma_data_HLC,
	dec_ma_data_DE, dec_ma_data_DEop1, dec_ma_data_DEop2,
	dec_ma_data_SPop1,
	dec_ma_data_BCop12, dec_ma_data_Bop12, dec_ma_data_Cop12,
	dec_sp_set_enable, dec_cpurd_enable, dec_cpuwr_enable,
	dec_mem_stage_op2, dec_mem_stage_op3, dec_mem_stage_op23,
	dec_prefix,
	stage_cut, A, X, B, C, D, E, H, L, CS, ES,
	buf2, buf1, buf0, ma, ma_pre, exma, maw1, slmem, slflash, slreg, slmirr, slexm, slbmem, sliram,
	imdr, cpuwr, cpuwr_reg, cpurd,
	hltst, stbst, dmama, dmarq, dmaack, waitdma, waitint, waitfl, waitexm, waitmod, waitmem, vcout,
	MAA, IE, SP, sp_inc, wdop, intdbg, intnmi, intrq3, intrq2, intrq1, intrq0,
	isp, intack, ivack, ivack_pre, monmd, monmdstp, softbrk, intisp,
	intblock, PSW_block, skp_block, wait_block_brtf,
	stage_cut_br, pc_set_brk, pc_set_dbg,
	prefix_ack, fchiram, fchiram_skp, romrd_skp, rstvec,
	flsize, bfsize, ramsize, bmsize, wait2nd,
	exmmsk, flmask, /*decdycut,*/ brkmsk,
	flread, fchram, mem_access,
// for EVA
        svi, svvcout,
        svintack, svmod, svmodf, svmodi,
        dec_alt1, dec_alt2, alt1, alt2,
        dec_sp_inc, idpop,
        flreadb,
        ID_stage3, ID_stage2,
        prefix, pcwaitf,
        icemsknmi, icemskdbg,
        cpumisal, sprel,
        pswen,
        // Ver1.51
        ocdmod,
//
	cpuen, baseck, resb, scanmode,
	dfsize, dflen,
	sldfwait_pre, sldflash, drdclk, waitdflash,
	wed, flspm, gofirm,
	RVEON, 
	gatead1, gatead2, gatead3, mdw,
	monpc, monma, monmdr, monmdw
	);

	output	[7:0]	ID_stage1, ID_stage0, ID_stage1_dec;
	output	[7:0]	MEM_stage1, MEM_stage0;
	output	[1:0]	stage_adr;
	output	[19:0]	pc, pc_inc;
	output		pc_wait_flg, stby_wait_flg, reg_wait, pa_data_buf, pa_data_mem;
	output		pa_data_spen;
	output		pa_st2;
	output	[17:0]	pa;
	output	[15:0]	ma, ma_pre;
	output	[3:0]	exma;
	output		maw1;
	output		slmem, slflash, slreg, slmirr, slexm, slbmem, sliram;
	output		intack, ivack, ivack_pre;
	output		monmd, monmdstp, softbrk;
	output		pc_set_brk, pc_set_dbg;
	output		prefix_ack, fchiram, fchiram_skp, romrd_skp;
	output		rstvec;
	output	[1:0]	intisp;
	output		data_hazard_flg, data_hazard, sp_hazard;
	output		INT_wait, wait2ndsfr, sl2ndwait_pre;
	output		dopen;
	output		brkmsk;
	output		flread, fchram;
	output		SP_enable, CS_enable;
	output		sldfwait_pre;
	output		sldflash;
	output		drdclk;
	output	[19:0]	monpc;
	output	[15:0]	monma;
	output	[15:0]	monmdr;
	output	[15:0]	monmdw;
// for EVA
        output          svintack, svmod, svmodf, svmodi;
        output          alt1, alt2;
        output          idpop;
        output  [3:0]   flreadb;
        output  [7:0]   ID_stage3, ID_stage2;
        output          prefix, pcwaitf;
        output          cpumisal;
        output          sprel;
	output		waitdflash;
//

	input	[31:0]	pid;
	input		dec_NMIS_enable;
	input		A_access,X_access,B_access,C_access;
	input		D_access,E_access,H_access,L_access;
	input		dec_RBS_enable, INT_access;
	input		dec_SP_enable;
	input		dec_pc_inc1, dec_pc_inc2, dec_pc_inc3, dec_pc_inc4, dec_clear_stage;
	input		dec_pc_set_enable;
	input		dec_pc_set_op01, dec_pc_set_op12, dec_pc_set_op123;
	input		dec_pc_set_AX, dec_pc_set_BC, dec_pc_set_DE, dec_pc_set_HL;
	input		dec_pc_set_pc1, dec_pc_set_pc2, dec_pc_set_pc3, dec_pc_set_pc12;
	input		dec_pc_set_calt, dec_pc_set_vec;
	input		dec_pc_set_brk, dec_pc_set_dbg;
	input		dec_pc_set_ret;
	input		dec_ma_enable;
	input		dec_ma_data_sp;
	input		dec_ma_data_saddr_op1, dec_ma_data_saddr_op2;
	input		dec_ma_data_sfr_op1, dec_ma_data_sfr_op2;
	input		dec_ma_data_op12, dec_ma_data_op23;
	input		dec_ma_data_HL, dec_ma_data_HLop1, dec_ma_data_HLop2;
	input		dec_ma_data_HLB, dec_ma_data_HLC;
	input		dec_ma_data_SPop1;
	input		dec_ma_data_DE, dec_ma_data_DEop1, dec_ma_data_DEop2;
	input		dec_ma_data_BCop12, dec_ma_data_Bop12, dec_ma_data_Cop12;
	input		dec_sp_set_enable;
	input		dec_cpurd_enable, dec_cpuwr_enable;
	input		dec_mem_stage_op2, dec_mem_stage_op3, dec_mem_stage_op23;
	input		dec_prefix;
	input		stage_cut;
	input	[7:0]	A, X, B, C, D, E, H, L, buf1, buf0;
	input		MAA;
	input	[3:0]	CS, ES, buf2;
	input	[15:0]	imdr;
	input	[15:0]	dmama;
	input		dmarq, dmaack, waitdma, waitint, waitfl, waitexm, waitmod, waitmem;
	input		hltst;
	input		stbst;		// add v1.50 2007.07.02 K.Tanaka
	input	[5:0]	vcout;
	input		IE;
	input	[14:0]	SP, sp_inc;
	input		wdop;
	input	[1:0]	isp;
	input		intdbg, intnmi, intrq3, intrq2, intrq1, intrq0;
	input		intblock, PSW_block, skp_block;
	input		wait_block_brtf;
	input		stage_cut_br;
	input	[3:0]	flsize, bfsize;
	input	[7:0]	ramsize;
	input	[3:0]	bmsize;
	input	[7:0]	wait2nd;
	input		cpuwr, cpuwr_reg, cpurd;
	input		exmmsk;
	input		flmask;
//	input		decdycut;
	input		mem_access;
	input		cpuen, baseck, resb;
	input		scanmode;
	input	[1:0]	dfsize;
	input		wed;
	input		flspm;
	input		gofirm;
	input		RVEON;
	input		gatead1, gatead2, gatead3;
	input	[15:0]	mdw;
// for EVA
        input           svi;
        input   [7:0]   svvcout;
        input           dec_alt1, dec_alt2;
        input           dec_sp_inc;
        input           icemsknmi, icemskdbg;
        input           pswen;
        input           ocdmod;
	input		dflen;
//

	wire	[15:0]	ma;
	wire	[3:0]	DS;
	wire	[17:0]	pa;
	wire	[1:0]	distance_pa_pc, pa_inc_en;
	wire		pa_st0, pa_st1, pa_st2, pa_st3;
	wire		pc_jump_en, pc_jump, pa_jump_en;
	wire		inc_pa;
	wire		pc_wait_flg, stby_wait_flg;
	wire	[18:0]	adrg, adrp;
	wire		adrsp1, adrsp2, adrsp3, adrsg0, adrsg1, adrsg2, adrsg3;
	wire		adrcy1, adrcy2, adrcy3, adrcy4;
	wire	[3:0]	adrout1, adrout2, adrout3, adrout4, adrout5;
	wire	[19:0]	adrout_ma, adrout_pa;
	wire		fchiram_wait, fchiram_ramrd, fchiram_romrd, prefix_wait;
	wire		pa_data_en, pa_data_sub2, pa_data_sub4;
	wire		brunch_en;
	wire		slexm_pre, slexm_pre2;
	wire		slram, slflash, slexm;
	wire		slmem_msk;
	wire		ma_data_saddr_op1a, ma_data_saddr_op1b, ma_data_saddr_op2a, ma_data_saddr_op2b;
	wire		ma_data_adrout, pc_set_adrout;
	wire		sp_hazard_flg, data_hazard_flg;
	wire		iopen, inten, nmien;
	wire		mirror_en, slmirr;
	wire		int_suspend, nmi_suspend, dma_suspend;
	wire		data_hazard_flg_pre;
	wire		pc_set_rp;
	wire		prefix_exe;
	wire		check234map_13, check234map_12, check234map_11, check234map_10;
	wire		check234map_03, check234map_02, check234map_01;
	wire		intclk_on;
	wire		SP_enable, CS_enable;
	wire	[15:0]	imdr_groupC;
	wire		sl2ndwait_pre, sl2ndwait_0, sl2ndwait_1, sl2ndwait_2, sl2ndwait_3, sl2ndwait_4, sl2ndwait_5, sl2ndwait_6, sl2ndwait_7, sl2ndwait;
	wire		dflash_countend_b;
//	wire		sldfwait_pre;
	wire		sldfwait;
	wire		intack_internal;
	wire		gatead;

	reg	[7:0]	ID_stage3, ID_stage2, ID_stage1, ID_stage0, ID_stage1_dec;
	reg	[7:0]	MEM_stage1, MEM_stage0;
	reg	[1:0]	stage_adr;
	reg	[19:0]	pc, pc_jump_address;
	reg	[19:0]	maw;
	reg	[15:0]	ma_pre;
	reg	[3:0]	exma;
	reg		slmem_pre, slreg, slexm_en, slflash_pre;
	reg		ma_enable_fchiram;
	reg	[17:0]	pa_pre;
	reg	[31:0]	id_que1;
	reg		inc_pa_pre, inc_pa_mst, inc_pa_slv;
	reg	[1:0]	pc_wait_cnt;
	reg		pc_wait_slv;
	reg		fchiram_wait_pre;
	reg		romrd_wait;
	reg		inc_que_flg;
	reg	[19:0]	pc_inc;
	reg		intack_pre, ivack_pre, ivack_end, ivack;
	reg		fchiram_pre;
	reg		ma_enable_slv;
	reg		prefix_ack, prefix_es;
	reg		pc_set_op01 ;
	reg		pc_set_brk, pc_set_dbg ;
	reg		pa_data_pre, pa_data_maw, pa_data_buf, pa_data_mem, pa_data_block;
	reg		pa_data_mlt1, pa_data_cyc1;
	reg	[19:0]	adrin1_ma, adrin1_pa, adrin2_ma, adrin2_pa, adrout_sub;
	reg		data_hazard, sp_hazard;
	reg		mkiack;
	reg		nmiack_buf, mkiack_buf;
	reg	[1:0]	intisp, intisp_pre;
	reg		int_suspend_fchiram;
	reg		inten_block, nmien_block;
	reg	[5:0]	vcode;
	reg		nmiack, dbgd, nmid, DBGS, NMIS;
	reg		monmd_pre, monmdstp_pre;
	reg		hazard_dbgintack;
	reg		softbrk;
	reg		rstvec;
	reg		SP_enable_pre, CS_enable_pre;
	reg		wait2ndsfr;
	reg		sldflash_enable;
	reg	[1:0]	dflash_count;
	reg		waitdflash;
	reg		sldflash;
	reg		drdclk;
	reg	[19:0]	pc_set_op01_data;

// for EVA
        reg             alt1i;
        reg             sviack, svintack, sviack_buf;
//

/*------------------------------------------------------------------------------*/
/* ���ɥ쥹�׻�(�����ѥ��ɥ쥹�׻�)                                           */
/*------------------------------------------------------------------------------*/
/* Ver2.0�������ѥ��ɥ쥹�黻���ʬ��						*/
/*------------------------------------------------------------------------------*/
// ���ɥ쥹�׻������ϣ�������
// ����դ�ʬ��̿��Ǥ��ä���硢�������Ω���ϡ�pa_pre���ɤߤ�����

	always @(dec_ma_data_BCop12 or dec_ma_data_DEop1 or dec_ma_data_DEop2 or
		dec_ma_data_HLop1 or dec_ma_data_HLop2 or dec_ma_data_HLB or dec_ma_data_HLC or
		dec_ma_data_SPop1 or dec_ma_data_Bop12 or dec_ma_data_Cop12 or
		B or C or D or E or H or L or DS or SP) begin
		case(1'b1)
			dec_ma_data_BCop12      : adrin1_ma = {DS,B,C} ;
			dec_ma_data_DEop1       : adrin1_ma = {DS,D,E} ;
			dec_ma_data_DEop2       : adrin1_ma = {DS,D,E} ;
			dec_ma_data_HLop1       : adrin1_ma = {DS,H,L} ;
			dec_ma_data_HLop2       : adrin1_ma = {DS,H,L} ;
			dec_ma_data_HLB         : adrin1_ma = {DS,H,L} ;
			dec_ma_data_HLC         : adrin1_ma = {DS,H,L} ;
			dec_ma_data_SPop1       : adrin1_ma = {4'hf,SP,1'b0} ;
			dec_ma_data_Bop12       : adrin1_ma = {DS,8'h00,B} ;
			dec_ma_data_Cop12       : adrin1_ma = {DS,8'h00,C} ;
			default                 : adrin1_ma = 20'h00000 ;
		endcase
	end

// ���ɥ쥹�׻������ϣ�������
	always @(dec_ma_data_HLop1 or dec_ma_data_DEop1 or dec_ma_data_SPop1 or
		dec_ma_data_HLop2 or dec_ma_data_DEop2 or
		dec_ma_data_BCop12 or dec_ma_data_Bop12 or dec_ma_data_Cop12 or
		dec_ma_data_HLB or dec_ma_data_HLC or
		ID_stage1 or ID_stage2 or B or C) begin
		case(1'b1)
			dec_ma_data_HLop1       : adrin2_ma = {12'h000,ID_stage1} ;
			dec_ma_data_DEop1       : adrin2_ma = {12'h000,ID_stage1} ;
			dec_ma_data_SPop1       : adrin2_ma = {12'h000,ID_stage1} ;
			dec_ma_data_HLop2       : adrin2_ma = {12'h000,ID_stage2} ;
			dec_ma_data_DEop2       : adrin2_ma = {12'h000,ID_stage2} ;
			dec_ma_data_BCop12      : adrin2_ma = {4'h0,ID_stage2,ID_stage1} ;
			dec_ma_data_Bop12       : adrin2_ma = {4'h0,ID_stage2,ID_stage1} ;
			dec_ma_data_Cop12       : adrin2_ma = {4'h0,ID_stage2,ID_stage1} ;
			dec_ma_data_HLB         : adrin2_ma = {12'h000,B} ;
			dec_ma_data_HLC         : adrin2_ma = {12'h000,C} ;
			default                 : adrin2_ma = 20'h00000 ;
		endcase
	end

// ���ɥ쥹�׻�

        assign adrout_ma = adrin1_ma + adrin2_ma;

/*------------------------------------------------------------------------------*/
/* ���ɥ쥹�׻�(���ʬ���ѥ��ɥ쥹�׻���                                        */
/*------------------------------------------------------------------------------*/
/* Ver2.0���ץ�����ѥ��ɥ쥹�黻���ʬ��					*/
/*------------------------------------------------------------------------------*/

// ���ɥ쥹�׻������ϣ�������
// ����դ�ʬ��̿��Ǥ��ä���硢�������Ω���ϡ�pa_pre���ɤߤ�����
	always @(dec_pc_set_pc1 or dec_pc_set_pc2 or dec_pc_set_pc3 or dec_pc_set_pc12 or pc_inc) begin
		case(1'b1)
			dec_pc_set_pc1  : adrin1_pa = pc_inc ;
			dec_pc_set_pc2  : adrin1_pa = pc_inc ;
			dec_pc_set_pc3  : adrin1_pa = pc_inc ;
			dec_pc_set_pc12 : adrin1_pa = pc_inc ;
			default         : adrin1_pa = 20'h00000 ;
		endcase
	end

// ���ɥ쥹�׻������ϣ�������
// ʬ���������Ω��(stage_cut)�ˡ����פʥ��ɥ쥹�׻��򤵤��ʤ���
	always @(dec_pc_set_pc1 or dec_pc_set_pc2 or dec_pc_set_pc3 or dec_pc_set_pc12 or
		ID_stage1 or ID_stage2 or ID_stage3) begin
		case(1'b1)
			dec_pc_set_pc1	: adrin2_pa = {{12{ID_stage1[7]}},ID_stage1} ;
			dec_pc_set_pc2	: adrin2_pa = {{12{ID_stage2[7]}},ID_stage2} ;
			dec_pc_set_pc3	: adrin2_pa = {{12{ID_stage3[7]}},ID_stage3} ;
			dec_pc_set_pc12	: adrin2_pa = {{4{ID_stage2[7]}},ID_stage2,ID_stage1} ;
			default		: adrin2_pa = 20'h00000 ;
		endcase
	end

// ���ɥ쥹�׻�

        assign adrout_pa = (stage_cut) ? {pa_pre[17:0],2'b0} : (adrin1_pa + adrin2_pa);

/*------------------------------------------------------------------------------*/
/* ���ɥ쥹�׻�(RAM�ե��å����Υե��å����ɥ쥹��                               */
/*------------------------------------------------------------------------------*/
/* Ver2.0��RAM�ե��å��ѥ��ɥ쥹�黻���ʬ��					*/
/*------------------------------------------------------------------------------*/

// RAM�ե��å����档fchiram���PC�Υ�����ȥ��åפ�Ϣư������ma�⥫����ȥ��åפ��뤬��
// ̿������ɤߤ���ɬ�פ����뤿�ᡢPC�λؤ����ɥ쥹����-4���뤤��-2����ma�򹹿����롣
// �ʲ���-2�������-4������ξ�����Ū�ˤϸ�ߤ˸�������뤬��RAM���֤˥����פ���ľ��ʤɤ�-2��
// ʬ�����Υ��ɥ쥹�黻��ͥ�褵���Τǡ�ʬ��Ƚ����Ǥ⡢pa_data_en��ͭ���ˤ��Ƥ�����ʤ���
	assign pa_data_en = fchiram & ~(dec_ma_enable) ;
	assign pa_data_sub2 = pa_data_en & ((pc_wait_cnt[1] | pc_wait_cnt[0]) | (fchiram_wait & (pc_wait_cnt == 1))) ;
	assign pa_data_sub4 = pa_data_en & (pc_wait_cnt == 2'b0) ;

	always @(pa_data_sub2 or pa_data_sub4 or pa_pre) begin
		case(1'b1)
			pa_data_sub2	: adrout_sub = {pa_pre[17:0],2'b0} - 2 ;
			pa_data_sub4	: adrout_sub = {pa_pre[17:0],2'b0} - 4 ;
			default		: adrout_sub = 20'h00000 ;
		endcase
	end

/*------------------------------------------------------------------------------*/
/* ������̿��¹ԥե饰							*/
/*------------------------------------------------------------------------------*/
/*   ������꥿����ʬ��̿��ǥץ���५���󥿤�ʬ����¹Ԥ���ե饰��������	*/
/*   �ңϣͥǡ������������κݤϡ��ץ���ॢ�ɥ쥹�Τߤ����濮����������롣	*/
/*------------------------------------------------------------------------------*/

// �ޥ����������̿��ν�λ���˥����פμ¹Ե��Ŀ��档
// ���ʬ��̿��Ǿ������Ω�Ȥʤä����ϣ��ˤʤ�ʬ���μ¹Ԥ��ޤ��롣
	assign brunch_en = ((stage_adr == 1) || (stage_adr == 2)) & stage_cut ;

// �ץ���५���󥿤Υ����׾�
// �����׼¹Ե��ľ��֤ǥ�����̿�᤬�ǥ����ɤ��줿��磱�ˤʤ롣
	assign pc_jump = (pc_set_op01 | pc_set_adrout |
			 dec_pc_set_op12 | dec_pc_set_op123 |
			 dec_pc_set_AX | dec_pc_set_BC | dec_pc_set_DE | dec_pc_set_HL |
			 dec_pc_set_calt | dec_pc_set_vec | dec_pc_set_brk | dec_pc_set_dbg) & ~brunch_en ;

// �ץ���५���󥿤Υ����׵��Ŀ��档
// ������̿��μ¹ԡ��꥿����̿��μ¹Ԥǣ��ˤʤ롣
// FLASH�Υǡ����ˤ����ʬ���Ǿ������Ω�Ȥʤä����ϣ��ˤʤ롣
// SP�ι�����ʬ��̿���Hazard��ȯ���������ϡ�ʬ��ư���ȯ�������餻�뤿�ᣱ����å�ʬ���ˤʤ롣
	assign pc_jump_en = (pc_jump | dec_pc_set_ret) & ~(pa_data_mem & ~stage_cut) & ~sp_hazard_flg;

// �ץ���ॢ�ɥ쥹���Ե�§�Ѳ����Ŀ��档
// FLASH�˥ǡ���������������ݤ�PC��̵�뤷��PA��񤭴�����ݤˣ��ˤʤ롣
	assign pa_jump_en = (pa_st3 & (pa_data_maw | prefix_wait | slmirr)) | pa_data_buf | pa_data_mlt1 | pa_data_cyc1 ;

/*------------------------------------------------------------------------------*/
/* �������襢�ɥ쥹����							*/
/*------------------------------------------------------------------------------*/
/*   ���������̿�����(�ңϣ�)���ɥ쥹�����򤹤롣				*/
/*------------------------------------------------------------------------------*/

// �٥������ɥ쥹�μ����߿��档
// �����������Ȥ��ݻ�����٤˰��ټ���ľ����
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)			pc_set_op01 <= 1'b0 ;
		else if (cpuen) begin
			if (pc_wait_flg)	pc_set_op01 <= pc_set_op01 ;
			else			pc_set_op01 <= dec_pc_set_op01 ;
		end
	end

// ���եȥ������֥졼�����档
// �����������Ȥ��ݻ�����٤˰��ټ���ľ����
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)			pc_set_brk <= 1'b0 ;
		else if (cpuen) begin
			if (pc_wait_flg)	pc_set_brk <= pc_set_brk ;
			else			pc_set_brk <= dec_pc_set_brk ;
		end
	end

// �ǥХå������߿��档
// �����������Ȥ��ݻ�����٤˰��ټ���ľ����
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)			pc_set_dbg <= 1'b0 ;
		else if (cpuen) begin
			if (pc_wait_flg)	pc_set_dbg <= pc_set_dbg ;
			else			pc_set_dbg <= dec_pc_set_dbg ;
		end
	end

// �٥��������ɤμ����ߡ�
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)			vcode <= 6'b0 ;
		else if (cpuen) begin
			if (data_hazard)	vcode <= vcode ;
// for EVA
                        else if (svintack | svmod | svmodi)     vcode <= svvcout[6:1] ;
//
			else			vcode <= vcout ;
		end
	end

// PC���Ф�ʬ��̿��ǥ��ɥ쥹�׻�����Ϥ����򤹤��
	assign pc_set_adrout = dec_pc_set_pc1 | dec_pc_set_pc2 | dec_pc_set_pc3 | dec_pc_set_pc12 ;

// ��������Υץ���५�����ͤ���˱��������ꡣ
/*------------------------------------------------------------------------------*/
/* Ver2.0��caseʸ���ѹ���SLFLASH�Υ��ԡ��ɥ��åפ򤷤䤹�������		*/
/*���������黻���adrout��ץ���ॢ�ɥ쥹�Ѥ�adrout_pa���ѹ�			*/
/*------------------------------------------------------------------------------*/
	always @(adrout_pa or
		 pc_set_op01 or dec_pc_set_op12 or dec_pc_set_op123 or pc_set_adrout or
		 dec_pc_set_AX or dec_pc_set_BC or dec_pc_set_DE or dec_pc_set_HL or
		 dec_pc_set_calt or dec_pc_set_vec or dec_pc_set_brk or dec_pc_set_dbg or
		 dec_pc_set_ret or pc or
		 ID_stage1 or ID_stage2 or ID_stage3 or vcode or
		 A or X or B or C or D or E or H or L or CS or
		 buf2 or buf1 or buf0 or pc_set_op01_data) begin
                case(1'b1)
                        pc_set_adrout           : pc_jump_address = adrout_pa ;
//                      pc_set_op01             : pc_jump_address = {4'b0, ID_stage3, ID_stage2} ;
			pc_set_op01             : pc_jump_address = pc_set_op01_data ;
                        dec_pc_set_op12         : pc_jump_address = {4'h0, ID_stage2, ID_stage1} ;
                        dec_pc_set_op123        : pc_jump_address = {ID_stage3[3:0], ID_stage2, ID_stage1} ;
                        dec_pc_set_AX           : pc_jump_address = {CS, A, X} ;
                        dec_pc_set_BC           : pc_jump_address = {CS, B, C} ;
                        dec_pc_set_DE           : pc_jump_address = {CS, D, E} ;
                        dec_pc_set_HL           : pc_jump_address = {CS, H, L} ;
                        dec_pc_set_calt         : pc_jump_address = {4'b0, 8'h00, 2'b10, ID_stage1[1:0], ID_stage1[6:4], 1'b0} ;
                        dec_pc_set_vec          : pc_jump_address = {4'b0, 8'h00, 1'b0, vcode, 1'b0} ;
                        dec_pc_set_brk          : pc_jump_address = {4'b0, 8'h00, 8'h7e} ;
                        dec_pc_set_dbg          : pc_jump_address = {4'b0, 8'h00, 8'h02} ;
                        dec_pc_set_ret          : pc_jump_address = {buf2, buf1, buf0} ;
                        default                 : pc_jump_address = pc ;
                endcase
	end

/*------------------------------------------------------------------------------*/
/* Ver3.0 ������ȯ�����Υ���������ѹ�					*/
/*��������pc_set_op01�λ���ʬ�����⡼��������				*/
/*------------------------------------------------------------------------------*/
	always @(svmod or pc or gofirm or monmd or ivack or flspm or RVEON or wed or ID_stage2 or ID_stage3) begin
		if (!svmod) begin
			if(pc == 20'h0 & gofirm) 	pc_set_op01_data <= 20'hEFFFC ;
			else if (monmd) begin
				if(flspm)	pc_set_op01_data <= 20'hF07E0 ;
				else 		pc_set_op01_data <= 20'hEFFF4 ;
			end
			else if(RVEON & ~wed & ivack)	pc_set_op01_data <= 20'hF08C0 ;
			else			pc_set_op01_data <= {4'h0, ID_stage3, ID_stage2} ;
		end
		else		pc_set_op01_data <= {4'h0, ID_stage3, ID_stage2} ;
	end
/*------------------------------------------------------------------------------*/
/* �ǡ�������(�ң���)�����̿��ե��å�����					*/
/*------------------------------------------------------------------------------*/
/*   �ץ���५���󥿤��ң��ͥ��ɥ쥹��ؤ��Ƥ����硢�ң��ͥե��å��⡼��	*/
/*   �����롣�������ңϣͥǡ������������κݤˤϡ����Υ⡼�ɤ���ȴ���롣		*/
/*------------------------------------------------------------------------------*/

// PC��RAM���֤�ؤ����ϡ��ʲ��ο��椬���ˤʤ�RAM�ե��å��򳫻Ϥ��롣
// FLASH�Υǡ����꡼�ɤȳ����߽����μ¹Ի��ˤϣ��ˤʤ롣
// FLASH�꡼�ɤ�fchiram�������Ȥ��Τϡ�FLASH���ɤ߽Ф���������Τߡ�
	assign fchiram = fchiram_pre & ~(pa_data_maw | pa_data_buf | pa_data_mlt1 | ivack) ;

// RAM���֤ؤΥե��å����������򼨤����档�ǡ������������ξ��ϣ��ˤʤ롣
// for EVA
//	assign fchram = fchiram & ~mem_access ;
        assign fchram = ((fchiram & ~mem_access) | (fchiram_pre & svintack)) ;
//

// PC��RAM���֤�ؤ��Ƥ��ʤ���硢�����פ����硢
// ES��Ȥä��ǡ������������ǥ��ɥ쥹��FLASH���֤�ؤ��Ƥ��ʤ��ä����˼��Υ���å���fchiram�򣰤ˤ��롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)		fchiram_pre <= 1'b0 ;
		else if (cpuen) begin
			if (pc_wait_flg)	fchiram_pre <= fchiram_pre ;
			else if (((pc_jump_address[19:16] > flsize) & (pc_jump_address[19:10] < {4'hE,2'b11,bfsize})) ||
				 (pc_jump_address[19:16] == 4'hf)) begin
				if (dec_sp_set_enable && pa_st3 && pc_jump_en)
						fchiram_pre <= 1'b0 ;
				else		fchiram_pre <= 1'b1 ;
			end
			else	fchiram_pre <= 1'b0 ;
		end
	end

/*------------------------------------------------------------------------------*/
/* �ңϣͥǡ���������������							*/
/*------------------------------------------------------------------------------*/
/*   �ߥ顼���֤�ţӤ�Ȥäƣңϣͤ˥ǡ���������������̿�᤬�¹Ԥ��줿��硢	*/
/*   �ѥ��ץ饤��������Ф���̿��Х�����ǡ������ɤ߽Ф������κݡ��¹�	*/
/*   ����������˱��������濮����������������롣				*/
/*------------------------------------------------------------------------------*/

// �ߥ顼���֥����������Ŀ��档ma���ߥ顼���֤���ꤷ����磱�ˤʤ롣
// for EVA
//	assign mirror_en = (maw[19:9] >= {4'hF,3'b000,bmsize}) & (maw[19:8] < {4'hf,ramsize}) ;
        assign mirror_en = (((svmodi || svmod) && !alt1i) ? 1'b0 : ((maw[19:9] >= {4'hF,3'b000,bmsize}) & (maw[19:8] < {4'hf,ramsize}))) & ~sldfwait_pre ;
//

// �ߥ顼�������򿮹档
// FLASH�Υǡ����꡼��ľ�塢�ޥ����������Ǥ�FLASH�ǡ��������������ϣ��ˤʤ롣
// FLASH�꡼�ɸ�ˡ�slmirr����Ȥ������~pa_data_mem��~pa_data_mlt1����Ѥ��롣
	assign slmirr = dec_cpurd_enable & mirror_en & ~pa_data_mem & ~pa_data_mlt1 ;

// RAM�������򿮹档
// �ߥ顼����������ˤϣ��ˤʤ롣
	assign slram = ~slmirr & (maw[19:16] == 4'hf) ;

// ����RAM�����򤵤줿�����Ȥʤ롣
	assign sliram = (
			 (( maw[15:9] < {3'b000,bmsize} ) |
			  ((maw[15:4] < {12'hFEE}) & (maw[15:8] >= {ramsize}))) &
			 ( maw[19:16] == 4'hf )) |
			(dmaack | exmmsk) ;

// for EVA

        reg             prefix;

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb)                              prefix <= 1'b0 ;
                else if (cpuen) begin
                        if (pc_wait_flg)                prefix <= prefix ;
                        else if (pa_st2)                prefix <= 1'b0 ;
                        else if (pa_data_maw)           prefix <= prefix ;
                        else if (pa_data_buf)           prefix <= prefix ;
                        else if (!dec_clear_stage)      prefix <= prefix ;
                        else if (prefix_ack && fchiram && dec_ma_enable)
                                                        prefix <= prefix ;
                        else                            prefix <= dec_prefix ;
                end
        end

        wire            prefix_block;

        assign prefix_block = (ID_stage0 == 8'hFF) | ({ID_stage0,ID_stage1} == 16'h61A1) |
                                 ({ID_stage0,ID_stage1} == 16'h61B1) | ({ID_stage0,ID_stage1} == 16'h61C1) ;
//

// FLASH�ؤΥǡ�����������ȯ����ɽ�����档
// �ǡ����ϥ����ɤ�ȯ���������ʳ��Υߥ顼���֥������������PREFIX̿��¹Ի��ˣ��ˤʤꡢ
// FLASH�ؤΥǡ���������������ݻ�����롣FLASH�꡼�ɥ�������ľ��ϣ��ˤʤ롣
// �ޥ����������̿��Σ�����å��ܤǤ�prefix_ack��Ω���夲��ESϢư��ͭ���ˤ��롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)				prefix_ack <= 1'b0 ;
		else if (cpuen) begin
			if (pc_wait_flg)			prefix_ack <= prefix_ack ;
			else if (slmirr && !data_hazard_flg)	prefix_ack <= 1'b1 ;
			else if (pa_st2)			prefix_ack <= 1'b0 ;
			else if (!dec_clear_stage && (stage_adr == 2'b00))
								prefix_ack <= prefix_ack ;
			else if (pa_data_maw)			prefix_ack <= prefix_ack ;
			else if (pa_data_buf)			prefix_ack <= prefix_ack ;
			else					prefix_ack <= dec_prefix | slmirr ;
		end
	end

// ����������̿���EXMEM���������Ǥϥ��ɥ쥹��ES��Ϣư������֤��Ĺ���롣
// prefix_ack��̿�ᥭ�塼������˻��Ѥ��Ƥ��뤿�ᡢ���̤ο�����б����롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)			prefix_es <= 1'b0 ;
		else if (cpuen) begin
			if (pc_wait_flg)	prefix_es <= prefix_es ;
			else if (!dec_clear_stage && (stage_adr == 2'b01))
						prefix_es <= prefix_ack ;
			else			prefix_es <= 1'b0 ;
		end
	end

// PREFIX̿���ES��FLASH���ְʳ���ؤ��������̾�ư��򤹤롣
// FLASH���֤�ؤ������Ϥ��ο��椬���ȤʤꡢFLASH�꡼��ư��򤹤롣
	assign prefix_exe = (pa_data_sub2 | pa_data_sub4) ?
	     prefix_ack & (((adrout_sub[19:16] != 4'hf) & ((adrout_sub[19:16] <= flsize) | (adrout_sub[19:10] >= {4'hE,2'b11,bfsize}))) | pa_st2 ) :
	     prefix_ack & (((maw[19:16] != 4'hf) & ((maw[19:16] <= flsize) | (maw[19:10] >= {4'hE,2'b11,bfsize}))) | pa_st2 ) ;

// PREFIX̿��ˤ��FLASH�꡼�ɥ����������濮�档
// PREFIX̿��¹Ը�ˣ��ˤʤꡢFLASH�꡼�ɥ�������ľ��ϣ��ˤʤ롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)				pa_data_pre <= 1'b0 ;
		else if (cpuen) begin
			if (pc_wait_flg && dec_prefix)	pa_data_pre <= pa_data_pre ;
			else if (pa_st2)		pa_data_pre <= 1'b0 ;
			else				pa_data_pre <= dec_prefix ;
		end
	end

// PREFIX̿�ᤪ��ӥߥ顼���֥꡼�ɥ������������濮�档
// PREFIX̿�᤬�¹Ԥ��줿���ȥߥ顼���֤����򤵤줿���ˣ��Ȥʤ롣
// �ǡ����ϥ����ɤ�ȯ����������PREFIX̿���RAM���֤˥��������������ϣ��ˤʤ롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)				pa_data_maw <= 1'b0 ;
		else if (cpuen) begin
// for EVA
//			if (slram | slexm_pre | pa_data_maw | pa_data_buf | data_hazard_flg)
                        if (slram | slexm_pre | pa_data_maw | pa_data_buf | data_hazard_flg | prefix_block)
//
								pa_data_maw <= 1'b0 ;
			else if (pc_wait_flg && dec_prefix)	pa_data_maw <= pa_data_maw ;
			else					pa_data_maw <= pa_data_pre | slmirr ;
		end
	end

// PID�Х��Υǡ�����Хåե��˳�Ǽ�������濮�档
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)	pa_data_buf <= 1'b0 ;
		else if (cpuen) pa_data_buf <= pa_data_maw ;
	end

// FLASH�ؤΥǡ��������������ޥ����������̿��Ǽ¹Ԥ��줿����ɽ�����档
// FLASH�꡼�ɤΥޥ����������̿��Ǥ�����򼨤���
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)	pa_data_mlt1 <= 1'b0 ;
		else if (cpuen) begin
			if (!dec_clear_stage)	pa_data_mlt1 <= pa_data_buf | pa_data_mem ;
			else 			pa_data_mlt1 <= 1'b0 ;
		end
	end

// FLASH�ؤΥǡ�������������������å�̿��Ǽ¹Ԥ��줿����ɽ�����档
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)	pa_data_cyc1 <= 1'b0 ;
		else if (cpuen) begin
			if (!dec_clear_stage) pa_data_cyc1 <= pa_data_mlt1 ;
			else pa_data_cyc1 <= 1'b0 ;
		end
	end

// �Хåե��˼������FLASH�Υǡ�������᤹���濮�档
// �ޥ����������̿��ˤ��FLASH�����������ä�����ʣ������å�Ω���夬�롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)	pa_data_mem <= 1'b0 ;
		else if (cpuen) begin
			if (pc_jump_en) pa_data_mem <= 1'b0 ;
			else  pa_data_mem <= pa_data_buf | (pa_data_mlt1 & dec_clear_stage) | pa_data_cyc1 ;
		end
	end

// FLASH�ؤΥ꡼�ɥ�������̿�Ὢλľ����Ω���夬�ꡢ�����߼����դ���֥�å����롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)	pa_data_block <= 1'b0 ;
		else if (cpuen) begin
			if (pa_data_block || (stage_adr != 2'b0)) pa_data_block <= 1'b0 ;
			else pa_data_block <= pa_data_mem ;
		end
	end

// FLASH�ؤΥǡ�������������������򼨤����档
	assign flread = pa_data_maw | pa_data_buf ;

// for EVA

        reg     [3:0]   flreadb;

        always @(flread or ma or wdop) begin
                if (flread) begin
                        casex ({wdop,ma[1:0]})
                                3'b0_00 : flreadb = 4'b0001 ;
                                3'b0_01 : flreadb = 4'b0010 ;
                                3'b0_10 : flreadb = 4'b0100 ;
                                3'b0_11 : flreadb = 4'b1000 ;
                                3'b1_00 : flreadb = 4'b0011 ;
                                3'b1_10 : flreadb = 4'b1100 ;
                                default : flreadb = 4'b0000 ;
                        endcase
                end
                else    flreadb = 4'b0000 ;
        end
//

// SP�ι������㳰Ū�˵�������ˡ�FLASH�Υǡ�����������ľ���ʬ���������򸡽Ф��롣
// ��������SP���̿��¹���Ǥ��ä����Ͼ嵭������̵���Ȥ��롣
	assign pa_data_spen = pa_data_block & ~SP_enable ;

// FLASH�ե��å����FLASH�إǡ�����������������磱�Ȥʤ롣
// ̿��¹Ԥ�NOP���֤������륹���å��װ���
	assign romrd_skp = pa_data_mem & ~pa_data_mlt1 ;

/*------------------------------------------------------------------------------*/
/* �ң��ͥ��ɥ쥹����								*/
/*------------------------------------------------------------------------------*/
/*   �ң��ͥ��ɥ쥹�����򤹤롣�Уңţƣɣ�̿��ľ��Ǥ���УţӤ�Ϣư���롣	*/
/*------------------------------------------------------------------------------*/

// ���̤��saddr����������ɽ�����档
	assign ma_data_saddr_op1a = dec_ma_data_saddr_op1 & (ID_stage1[7:5] == 3'b000) ;
	assign ma_data_saddr_op1b = dec_ma_data_saddr_op1 & ~(ID_stage1[7:5] == 3'b000) ;
	assign ma_data_saddr_op2a = dec_ma_data_saddr_op2 & (ID_stage2[7:5] == 3'b000) ;
	assign ma_data_saddr_op2b = dec_ma_data_saddr_op2 & ~(ID_stage2[7:5] == 3'b000) ;

// �ǡ����������ȡ�PREFIX̿��¹Ի��ˤ�ES���֤�����롣
// for EVA
//	assign DS = (prefix_ack || prefix_es) ? ES : 4'hf ;
        assign DS = ((prefix_ack || prefix_es) && ~prefix_block) ? ES : 4'hf ;
//

// ���ɥ쥹�׻�����Ϥ�ma�Ȥ������򤹤뿮�档
	assign ma_data_adrout = dec_ma_data_HLop1 | dec_ma_data_HLop2 |
				dec_ma_data_HLB | dec_ma_data_HLC |
				dec_ma_data_DEop1 | dec_ma_data_DEop2 | dec_ma_data_SPop1 |
				dec_ma_data_BCop12 | dec_ma_data_Bop12 | dec_ma_data_Cop12 ;

// ���ɥ쥹����˱��������ꤹ�롣
// Hazard��ȯ����������RAM�ե��å����SP�ι�����ʬ��̿���Hazard��ȯ���������ϡ�
// �����ʥ��ꥢ���������ɤ����ᣰ�ˤʤ롣���ξ��SLMEM�⣰�ˤʤ롣
/*------------------------------------------------------------------------------*/
/* Ver2.0��pa_data_sub2,sub4��RAM�ե��å����η�ϩ��ma_pre�˥����쥯�Ȥ���³����	*/
/*�����������ΰ٤�maw����Ϻ�����롣maw��SLFLASH�ξ�����ि�ᡢSLFLASH��	*/
/*�����������ԡ��ɥ��åפ�Ԥʤ���						*/
/*���������黻���adrout����ꥢ�ɥ쥹�Ѥ�adrout_ma���ѹ�			*/
/*------------------------------------------------------------------------------*/
	always @(adrout_ma or DS or ma or D or E or H or L or
		 ID_stage1 or ID_stage2 or ID_stage3 or
		 dec_ma_data_sfr_op1 or dec_ma_data_sfr_op2 or
		 ma_data_saddr_op1a or ma_data_saddr_op2a or ma_data_saddr_op1b or ma_data_saddr_op2b or
		 dec_ma_data_op12 or dec_ma_data_op23 or dec_ma_data_DE or dec_ma_data_HL or
		 dec_ma_data_sp or ma_data_adrout or pc_jump_en or
		 sp_inc or sp_hazard_flg or data_hazard_flg or fchiram) begin
		if (data_hazard_flg && ~(fchiram && pc_jump_en && ~sp_hazard_flg))
						maw = 20'h00000 ;
		else if (ma_data_adrout)	maw = adrout_ma ;
		else if (ma_data_saddr_op1a)	maw = {DS, 8'hff, ID_stage1} ;
		else if (ma_data_saddr_op1b)	maw = {DS, 8'hfe, ID_stage1} ;
		else if (ma_data_saddr_op2a)	maw = {DS, 8'hff, ID_stage2} ;
		else if (ma_data_saddr_op2b)	maw = {DS, 8'hfe, ID_stage2} ;
		else if (dec_ma_data_sfr_op1)	maw = {DS, 8'hff, ID_stage1} ;
		else if (dec_ma_data_sfr_op2)	maw = {DS, 8'hff, ID_stage2} ;
		else if (dec_ma_data_op12)	maw = {DS, ID_stage2, ID_stage1} ;
		else if (dec_ma_data_op23)	maw = {DS, ID_stage3, ID_stage2} ;
		else if (dec_ma_data_DE)	maw = {DS, D, E} ;
		else if (dec_ma_data_HL)	maw = {DS, H, L} ;
		else if (dec_ma_data_sp)	maw = {DS, sp_inc, 1'b0} ;
		else				maw = 20'h00000 ;
	end

// FLASH�ǡ����꡼�ɻ��˥Хåե��˼�����PID�Х��ξ��¦������¦�������򤹤뿮�档
	assign maw1 = maw[1] ;

// for EVA

        reg             sprel;

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb) begin
                        sprel <= 1'b0 ;
                end
                else if (cpuen) begin
                        if (reg_wait) begin
                                sprel <= sprel ;
                        end
                        else begin
                                sprel <= dec_ma_data_SPop1 ;
                        end
                end
        end
//

/*------------------------------------------------------------------------------*/
/* �ң��ͥ��ɥ쥹�쥸����							*/
/*------------------------------------------------------------------------------*/
/*   �ң��ͥ��ɥ쥹���Ǽ���롣���ɥ쥹��������֤Τɤ��ΰ��ؤ��Ƥ��뤫��	*/
/*   Ƚ�ꤹ�롣�ң��ͥե��å���ң��ͥǡ�������������ȯ���������ϡ�		*/
/*   �ѥ��ץ饤��������Ф����濮����������롣				*/
/*------------------------------------------------------------------------------*/

// FLASH�ؤΥե��å�����������ɽ�����档
// PA��FLASH���֤�ؤ��Ƥ��ơ����ĥ��󥯥���Ȥ�������ˤʤ롣
// RAM�ե��å���ʤ�FLASH�˥ե��å������������ʤ����ϣ��ˤʤ롣
// for EVA
        wire erea_flash = (svmodf & ~(alt1i & alt1)) ? (pa[17:14] != 4'hf) :
                                                        ((pa[17:14] <= flsize) || (pa[17:8] >= {4'hE,2'b11,bfsize}) && (pa[17:14] != 4'hf)) ;
//
// PA���ե�å�����֤�ؤ��Ƥ���������о�
// ���ġ��ץ�ե��å�����(~pa_st3)���ޤ���PA������(inc_pa)���ޤ���ʬ���¹Ի�(pc_jump_en)��
// �ޤ���FLASH�ǡ���������������SLFLASH�򹹿����롣
// ��������FLASH�ǡ�����������̿�᤬�ޥ����������̿����ä����ϡ��ݻ�����ɬ�פ����롣
/*------------------------------------------------------------------------------*/
/* Ver2.0��SLFLASH�Υ��ԡ��ɥ��åפΤ��ᡢ�ͥå��Ȥʤ�slmirr��prefix_wait�ο���	*/
/*���������η�ϩ���ڤ롣							*/
/*        slmirr��Flash�꡼�ɤΣ�ȯ�ܤ�Ω�����������礭���Τ��Ѳ����ԡ��ɤ��٤�	*/
/*����������ȯ�ܤΥǡ����ϸ������Ѥ��Ƥ��ʤ����ᡢ¾�ο�����ѹ����롣		*/
/*�������������pa_data_maw(��ȯ�ܡˡ�pa_data_buf(��ȯ��)����Ѥ��롣		*/
/*------------------------------------------------------------------------------*/
// for EVA
//	always @(pa or flsize or bfsize or pa_st3 or inc_pa or pc_jump_en or pa_data_maw or pa_data_buf) begin
        always @(erea_flash or pa_st3 or inc_pa or pc_jump_en or pa_data_maw or pa_data_buf) begin
//
// for EVA
//		if (((pa[17:14] <= flsize) || (pa[17:8] >= {4'hE,2'b11,bfsize}) && (pa[17:14] != 4'hf))) begin
                if (erea_flash) begin
//
//			slflash_pre = ~pa_st3 | inc_pa | pc_jump_en | slmirr | prefix_wait ;
			slflash_pre = ~pa_st3 | inc_pa | pc_jump_en | pa_data_maw | pa_data_buf ;
//
		end
		else begin
			slflash_pre = 1'b0 ;
		end
	end

// FLASH�꡼�ɤ��ޥ����������̿��Ǥ��ä����(pa_data_mlt1)�ϡ�SLFLASH�����Ω��������PID�ǡ������ݻ����롣
// ��������ʬ����(pc_jump_en)��ʬ������Τǡ��ݻ����ʤ���
	assign slflash = ((slflash_pre & ~(pa_data_mlt1 & ~pc_jump_en)) | (pc == 0)) & flmask ;

// ��������ؤΥե��å����ǡ��������������ǣ��Ȥʤ롣
	always @(fchiram or dec_cpurd_enable or dec_cpuwr_enable or pa_st2) begin
		if (fchiram) begin
			slexm_en = (dec_cpuwr_enable & ~pa_st2) | (dec_cpurd_enable | ~dec_cpuwr_enable | pa_st2) ;
		end
		else begin
			slexm_en = dec_cpuwr_enable | dec_cpurd_enable ;
		end
	end

// ��������������򿮹档FLSIZE����ˤ�����򤵤줿�ϰϤǣ��Ȥʤ롣
// DMAž����ϣ��ȤʤꡣDMA�ȳ����Х���������Ȥζ�����򤱤롣
/*------------------------------------------------------------------------------*/
/* Ver2.0��maw(�ǡ����꡼��)�η�ϩ��ꡢRAM�ե��å����α黻����̤ˤ�����	*/
/*�����������ΰ١���������ե��å�����adrout_sub����Ѥ��뤿�ᡢ�������򿮹�	*/
/*        ���ɲá�								*/
/*------------------------------------------------------------------------------*/
// for EVA
//	assign slexm_pre = slexm_en & ((maw[19:16] > flsize) &	
//                (maw[19:10] < {4'hE,2'b11,bfsize}) & (maw[19:16] != 4'hf)) & ~(exmmsk | dmaack) ;
//	assign slexm_pre2 = slexm_en & ((adrout_sub[19:16] > flsize) &
//		(adrout_sub[19:10] < {4'hE,2'b11,bfsize}) & (adrout_sub[19:16] != 4'hf)) & ~(exmmsk | dmaack) ;
//
// for EVA
        wire erea_exmem = (svmodf & ~(alt1)) ? 1'b0 : ((maw[19:16] > flsize) & 
                (maw[19:10] < {4'hE,2'b11,bfsize}) & (maw[19:16] != 4'hf)) ;
        wire erea_exmem2= (svmodf & ~(alt1)) ? 1'b0 : ((adrout_sub[19:16] > flsize) & 
                (adrout_sub[19:10] < {4'hE,2'b11,bfsize}) & (adrout_sub[19:16] != 4'hf)) ;
//        assign slexm_pre = slexm_en & erea_exmem & ~(exmmsk | dmaack | wait2ndsfr) ;
//        assign slexm_pre2 = slexm_en & erea_exmem2 & ~(exmmsk | dmaack | wait2ndsfr) ;
        assign slexm_pre = slexm_en & erea_exmem & ~(exmmsk | dmaack | wait2ndsfr | waitdflash) ;
        assign slexm_pre2 = slexm_en & erea_exmem2 & ~(exmmsk | dmaack | wait2ndsfr | waitdflash) ;
//
	assign slexm = (pa_data_sub2 | pa_data_sub4) ?
			slexm_pre2 & ~(dec_ma_enable & fchiram & pc_wait_flg) :
			slexm_pre & ~(dec_ma_enable & fchiram & pc_wait_flg) ;

// RAM���ɥ쥹�ȶ������򿮹档�����ߤ䥸����̿��Υϥ����ɤ�������������ȯ�����ˤ��ݻ�����롣
/*------------------------------------------------------------------------------*/
/* Ver2.0��SLFLASH�Υ��ԡ��ɥ��åפΤ��ᡢpa_data_sub2,pa_data_sub4(RAM�ե��å�)*/
/*���������κݤϥ��ɥ쥹�黻������Ѥ˻�����ľ��adrout_sub�����Ϥ���褦���ѹ���*/
/*        dec_ma_enable����ma_pre��maw���ͤ�����Ƥ��뤬���ϥ�����ȯ�����ˣ���	*/
/*���������ʤäƤ��ޤ���maw���ϥ�����ȯ�����ˣ��ˤ��Ƥ��뤬��ma_pre�ˤϥϥ�����	*/
/*�����������ν��������äƤ��ʤ�����Ǥ��롣������maw�Υϥ����ɾ��ȯ������Ʊ��	*/
/*��������������ma_pre���ͤ��Ѥ��ʤ��褦�ˤ��롣				*/
/*------------------------------------------------------------------------------*/
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) begin
			exma <= 4'h0 ;
			ma_pre <= 16'h0000 ;
			slmem_pre <= 1'b0 ;
			slreg <= 1'b0 ;
		end
		else if (cpuen) begin
			if ((dec_pc_set_ret && pc_wait_flg) ||
			    (dec_sp_set_enable && (pc_wait_slv && !(data_hazard || sp_hazard)))) begin
				exma <= exma ;
				ma_pre <= ma_pre ;
				slmem_pre <= slmem_pre ;
				slreg <= slreg ;
			end
			else if ((pa_data_sub2 || pa_data_sub4) & ~(pc_set_adrout & ~stage_cut)) begin
				exma <= adrout_sub[19:16] ;
				ma_pre <= adrout_sub[15:0] ;
				if ((adrout_sub[19:16] == 4'hf) & !mirror_en) slmem_pre <= 1'b1 ;
				else                                          slmem_pre <= 1'b0 ;
				slreg <= 1'b0 ;
			end
			else if (dec_ma_enable || fchiram) begin
				exma <= maw[19:16] ;
				if (data_hazard_flg && ~(fchiram && pc_jump_en && ~sp_hazard_flg)) ma_pre <= ma_pre;
				else ma_pre <= maw[15:0] ;
				if (maw[19:5] == 15'h7ff7) begin
					slmem_pre <= 1'b0 ;
					slreg <= 1'b1 ;
				end
				else if ((maw[19:16] == 4'hf) & !mirror_en) begin
					slmem_pre <= 1'b1 ;
					slreg <= 1'b0 ;
				end
				else begin
					slmem_pre <= 1'b0 ;
					slreg <= 1'b0 ;
				end
			end
		end
	end

// RAM�ե��å����RAM�������������ݻ����档
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)	ma_enable_fchiram <= 1'b0 ;
		else if (cpuen)	ma_enable_fchiram <= dec_ma_enable & fchiram ;
	end

// slmem�Υޥ�����¿�ť����������ɤ���
// ���������������򿮹�ϡ��쥸�������ϤǤʤ��ƤϤ����ʤ����ᡢpc_wait_cnt��Ȥ���
// RAM�ե��å����HALT/STOP�˰ܹԤ������ϡ�RAM�ؤΥե��å������������ɤ���
	assign slmem_msk = (ma_enable_fchiram & (pc_wait_cnt[1] | pc_wait_cnt[0])) | waitfl | stbst ;	// add stbst v1.50 2007.07.02 K.Tanaka

// RAM�������򿮹档CPUWR��CPURD�����λ���Ω�ġ�
// DMAž�����̵����SLMEM�򣱤ˤ��롣
	assign slmem = (slmem_pre & (cpuwr | cpurd) & ~(slmem_msk)) | waitdma ;

// �ºݤ˽��Ϥ����ma����ɥ����������Ϻǲ��̥ӥåȤ�������ˤʤ������ϤؤΥ���������ػߤ��롣
// DMAž������dmama����Ϥ��롣���λ��������ϤؤΥ�ɥ��������϶ػߡ�
	assign ma = (waitdma) ? (wdop) ? {dmama[15:1],1'b0} : dmama : 
				(wdop) ? {ma_pre[15:1],1'b0} : ma_pre ;

// for EVA
        wire            cpumisal;

	// for EVA Ver2.01 RAM�ե��å���ϥǡ������������Τߤ˸��ꤹ�롣
        // assign cpumisal = wdop & ma_pre[0] & (cpuwr | cpurd) ;
	assign cpumisal = (!fchiram) ?  wdop & ma_pre[0] & (cpuwr | cpurd) :
					wdop & ma_pre[0] & (cpuwr | cpurd) & ma_enable_fchiram ;
//

// RAM�ե��å����RAM�ؤΥǡ�������������ȯ��������硢
// �ʲ��ο����̿�ᥭ�塼���ѥ��ץ饤��쥸�����������Ԥʤ���
// RAM�ե��å����̾�ξ��ʬ����ʬ�����ʤ���硢���ν��������פ�����
// FLASH�ǡ����򻲾Ȥ������ϡ�PA���ɤ�ľ�������򣲥���å����Ǽ¸����롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)				ma_enable_slv <= 1'b0 ;
		else if (cpuen) begin
			if (pc_wait_flg)		ma_enable_slv <= ma_enable_slv ;
			else if (dec_clear_stage)	ma_enable_slv <= (dec_ma_enable & ~pc_jump_en) | pa_data_mlt1 ;
		end
	end

/*------------------------------------------------------------------------------*/
/* Ver2.0 2ndSFR��������ȯ������						*/
/*------------------------------------------------------------------------------*/
/*   NPB�ޥ������ܤ���ݤΥ�������ȯ���Τ��ᡢ2ndSFR�ؤΥ����������˥�������	*/
/*   ��ȯ�������롣								*/
/*     F0000-F00FF  WAIT2ND0=1�ǥ�������					*/
/*     F0100-F01FF  WAIT2ND1=1�ǥ�������					*/
/*     F0200-F02FF  WAIT2ND2=1�ǥ�������					*/
/*     F0300-F03FF  WAIT2ND3=1�ǥ�������					*/
/*     F0400-F04FF  WAIT2ND4=1�ǥ�������					*/
/*     F0500-F05FF  WAIT2ND5=1�ǥ�������					*/
/*     F0600-F06FF  WAIT2ND6=1�ǥ�������					*/
/*     F0700-F07FF  WAIT2ND7=1�ǥ�������					*/
/*										*/
/*  exmmsk����ˤ�waitexm�����äƤ��ʤ������ΰ٤�waitexm���ɲä���ɬ�פ��ꡣ	*/
/*------------------------------------------------------------------------------*/

	assign sl2ndwait_0 = (maw[10:8] == 3'b000) & wait2nd[0] ;
	assign sl2ndwait_1 = (maw[10:8] == 3'b001) & wait2nd[1] ;
	assign sl2ndwait_2 = (maw[10:8] == 3'b010) & wait2nd[2] ;
	assign sl2ndwait_3 = (maw[10:8] == 3'b011) & wait2nd[3] ;
	assign sl2ndwait_4 = (maw[10:8] == 3'b100) & wait2nd[4] ;
	assign sl2ndwait_5 = (maw[10:8] == 3'b101) & wait2nd[5] ;
	assign sl2ndwait_6 = (maw[10:8] == 3'b110) & wait2nd[6] ;
	assign sl2ndwait_7 = (maw[10:8] == 3'b111) & wait2nd[7] ;

	assign sl2ndwait_pre = slexm_en & (maw[19:12] == 8'hf0) & (maw[11] == 1'b0) &
		(sl2ndwait_0 | sl2ndwait_1 | sl2ndwait_2 | sl2ndwait_3 | sl2ndwait_4 | sl2ndwait_5 | sl2ndwait_6 | sl2ndwait_7);

	assign sl2ndwait = sl2ndwait_pre & ~(dec_ma_enable & fchiram & pc_wait_flg) & ~(exmmsk | waitexm | waitdflash);

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if      (!resb)      wait2ndsfr <= 1'b0 ;
		else if (wait2ndsfr) wait2ndsfr <= waitmem ;
		else if (sl2ndwait)  wait2ndsfr <= 1'b1 ;
		else                 wait2ndsfr <= 1'b0 ;
	end

/*------------------------------------------------------------------------------*/
/* Ver3.0 Data_Flash��������ȯ������						*/
/*------------------------------------------------------------------------------*/
/*   DataFlash������������1����å����������Ǥϥ��ԡ��ɥͥå��ˤ뤿�ᥦ������	*/
/*   �б���»ܡ�								*/
/*     none  :		      DFSIZE[1:0] = 2'h00;				*/
/*     4K    : F1000H-F1FFFH  DFSIZE[1:0] = 2'h01;				*/
/*     8K    : F1000H-F2FFFH  DFSIZE[1:0] = 2'h10;				*/
/*     16K   : F1000H-F4FFFH  DFSIZE[1:0] = 2'h11;				*/
/*  exmmsk����ˤ�waitexm�����äƤ��ʤ������ΰ٤�waitexm���ɲä���ɬ�פ��ꡣ	*/
/*------------------------------------------------------------------------------*/

	always @(dfsize[1:0] or maw[14:12]) begin
		casex ({dfsize[1:0], maw[14:12]})
			{2'b00,3'bxxx} : sldflash_enable = 1'b0;
			{2'b01,3'b001} : sldflash_enable = 1'b1; /* F1000H-F1FFFH */
			{2'b10,3'b001} : sldflash_enable = 1'b1; /* F1000H-F2FFFH */
			{2'b10,3'b010} : sldflash_enable = 1'b1; /* F1000H-F2FFFH */
			{2'b11,3'b001} : sldflash_enable = 1'b1; /* F1000H-F4FFFH */
			{2'b11,3'b010} : sldflash_enable = 1'b1; /* F1000H-F4FFFH */
			{2'b11,3'b011} : sldflash_enable = 1'b1; /* F1000H-F4FFFH */
			{2'b11,3'b100} : sldflash_enable = 1'b1; /* F1000H-F4FFFH */
			default : sldflash_enable = 1'b0;
		endcase
	end

	assign sldfwait_pre = slexm_en & (maw[19:16] == 4'hf) & (maw[15] == 1'b0) & sldflash_enable;

	assign sldfwait = sldfwait_pre & ~(dec_ma_enable & fchiram & pc_wait_flg) & ~(exmmsk | waitexm | wait2ndsfr);

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if      (!resb)      		waitdflash <= 1'b0 ;
		else begin
			if (waitdflash) 	waitdflash <= dflash_countend_b ;
			else if (sldfwait)   	waitdflash <= 1'b1 ;
			else                 	waitdflash <= 1'b0 ;
		end
	end

	always @(posedge baseck or negedge resb) begin
		if	(!resb)	     		dflash_count <= 2'b10 ;
		else begin
			if (waitdflash) begin
				if (dflash_count == 2'b00)
					dflash_count <= 2'b10 ;
				else	dflash_count <= dflash_count - 1'b1 ;
			end
			else		     	dflash_count <= 2'b10 ;
		end
	end

	assign	dflash_countend_b = dflash_count[1] | dflash_count[0] ;

/*------------------------------------------------------------------------------*/
/* Ver3.0 SLDFLASH : DataFlash������������					*/
/*------------------------------------------------------------------------------*/

	always @(posedge baseck or negedge resb) begin
		if	(!resb)		sldflash <= 1'b0 ;
		else if	(dflen) begin
			if 	(!sldflash)	sldflash <= sldfwait ;
			else begin
				if (sldfwait || waitdflash)	sldflash <= 1'b1 ;
				else				sldflash <= 1'b0 ;
			end
		end
		else		sldflash <= 1'b0 ;
	end

/*------------------------------------------------------------------------------*/
/* Ver3.0 DRDCLK : DataFlash������������					*/
/*------------------------------------------------------------------------------*/

	always @(posedge baseck or negedge resb) begin
		if (!resb)		drdclk <= 1'b1 ;
		else if (dflen) begin
			if (waitdflash) begin
				if (dflash_count == 2'b01)	drdclk <= 1'b1 ;
				else				drdclk <= 1'b0 ;
			end
			else		drdclk <= 1'b1 ;
		end
		else			drdclk <= 1'b1 ;
	end

/*------------------------------------------------------------------------------*/
/* Ver2.0 SP,CS�쥸����������������						*/
/*------------------------------------------------------------------------------*/
/*   SP,CS�쥸�����ϥϥ������װ����뤿�ᡢSLFLASH�ؤΥ����ߥ󥰥ͥå��ѥ���	*/
/*   �ʤ롣���Τ��ᡢMEM���ơ����ǤϤʤ���ADR���ơ����ǥǥ����ɤ�Ԥʤ���	*/
/*------------------------------------------------------------------------------*/
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) begin
			SP_enable_pre <= 1'b0 ;
			CS_enable_pre <= 1'b0 ;
		end
		else if (cpuen & dec_ma_enable) begin
			if (maw[19:1] == 19'h7fffc) SP_enable_pre <= 1'b1 ;	//SP���ɥ쥹��FFFF8,FFFF9
			else                        SP_enable_pre <= 1'b0 ;
			if (maw[19:0] == 20'hffffc) CS_enable_pre <= 1'b1 ;	//CS���ɥ쥹��FFFFC
			else                        CS_enable_pre <= 1'b0 ;
		end
	end
	assign SP_enable = dec_SP_enable | (cpuwr_reg & SP_enable_pre);
	assign CS_enable = cpuwr_reg & CS_enable_pre;

/*------------------------------------------------------------------------------*/
/* ����������������								*/
/*------------------------------------------------------------------------------*/
/*   �ϥ�����ȯ�������ң��ͤؤΥե��å��������������ңϣͥǡ���������������	*/
/*   �ģͣ�ȯ�����������������ȿ����ȯ�������롣				*/
/*   ��������ȯ���װ��μ���ˤ�äƥ������Ȼ��֤����椹�롣			*/
/*------------------------------------------------------------------------------*/

// RAM�ե��å����������������ȯ���װ���
// RAM�ե��å���ξ��ʬ����FLASH�꡼�ɤʤɤ����RAM����������ɽ�����档
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)				fchiram_wait_pre <= 1'b0 ;
		else if (cpuen) begin
			if (pc_wait_flg)		fchiram_wait_pre <= fchiram_wait_pre ;
			else if (((pa_inc_en == 2'h1) || ((dec_ma_enable || stage_cut_br) && (dec_clear_stage || stage_cut)))
				 && (pa_inc_en != 2'h0) && ~(pa_data_buf && !inc_pa))
							fchiram_wait_pre <= 1'b1 ;
			else 				fchiram_wait_pre <= 1'b0 ;
		end
	end

// RAM�ե��å���������������ȿ��档PC�β��̣��ӥåȤ�2'b11���ä����ǡ�
// �嵭�ξ����������Ƥ���������������Ȥ�ȯ�����롣�������Ȼ��֤ϣ�����å���
// fchiram_ramrd�ϡ����Х���̿��ȡ�PC�����夬2'b11�Υ��ɥ쥹��ʬ����������Ω�ġ�
// �������Ȥ���������RAM�ե��å����ΥХ���������Ԥʤ���
	assign fchiram_wait = fchiram & pc[1] & pc[0] & ~dec_ma_enable & (dec_pc_inc4 || pa_st2) ;

// RAM�ե��å���������������ȿ��椬RAM����������ȯ��������磱�Ȥʤ롣
	assign fchiram_ramrd = fchiram_wait & ma_enable_slv ;

// RAM�ե��å����FLASH�꡼�ɥ���������ȯ��������磱�Ȥʤ롣
	assign fchiram_romrd = fchiram & prefix_exe & ~inc_pa_mst ;

// FLASH�ؤΥ꡼�ɥ�����������ȯ�������������������װ����������Ȼ��֤ϣ�����å���
// for EVA
//	assign prefix_wait = prefix_ack & (pa_data_pre | pa_data_maw | pa_data_buf) & ~slram & ~slexm_pre ;
        assign prefix_wait = prefix_ack & (pa_data_pre | pa_data_maw | pa_data_buf) & ~slram & ~slexm_pre & ~prefix_block ;
//

// FLASH�ե��å����FLASH�ؤΥ꡼�ɥ����������ˣ��Ȥʤ롣
// ������������ȯ���װ��ǤϤʤ���PA�Υ��󥯥���Ȥ�̿�ᥭ�塼��ž�������椹�롣
// FLASH�ؤΥǡ���������������PID�ǡ������ľ����ȯ�����롣�̾盧�ο��椬���Ǥ�
// PID�ǡ����μ��ľ���ͤˣ�����å��Υ������Ȥ����롣��������FLASH��������̿��¹Ի��ˡ�
// PA�Υ��󥯥���Ȥ�̵�����ϡ�PID�ǡ������ľ���Υ������Ȥ����פ�����
// �¹ԥ���å������碌�뤿��˸Ĥο���ǥ������Ȥ��������롣�ü��������פ��륱������
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)				romrd_wait <= 1'b0 ;
		else if (cpuen) begin
			if (pc_wait_flg & fchiram)	romrd_wait <= romrd_wait ;
			else if (~fchiram & (pa_data_buf || pa_data_mlt1 || pa_data_cyc1) & ~inc_pa)
							romrd_wait <= 1'b1 ;
			else 				romrd_wait <= 1'b0 ;
		end
	end

// �ºݤ������������ȿ��档�ǡ����ϥ�����ȯ�����Ϥ��ʤ餺���ˤʤ롣
// ����¾���װ���������������ľ��Ǥʤ����ˣ��Ȥʤ롣
	assign pc_wait_flg = (((fchiram & ~pa_st0) | prefix_wait | (slmirr & ~pa_data_mlt1)) & ~pc_wait_slv) | data_hazard_flg ;

/*------------------------------------------------------------------------------*/
/* Ver2.0 stby�ο��椬SLFLASH����ߥ��ԡ��ɥͥå��Ȥʤ뤿�ᡢ�ϥ����ɾ���	*/
/*��������ȴ����stby_wait_flg�������						*/
/*------------------------------------------------------------------------------*/
	assign stby_wait_flg = fchiram & ~pa_st0 & ~pc_wait_slv ;

// ������ư���INT�ޥ����IF/MK�쥸������PSW�ؤΥ饤�ȥ������������礹��������ꤷ��
// �����������Ȥ�ȯ�������롣������RETI/RETB̿�ᡢ�����������ȤǤ�ȯ�����ʤ���
	assign INT_wait = (INT_access | (slmem_pre & cpuwr & ((ma[15:0] == 16'hfffa) | (ma[15:4] == 12'hffe) | (ma[15:4] == 12'hffd))))
			 & ~({ID_stage0,ID_stage1} == 16'h61FC) & ~({ID_stage0,ID_stage1} == 16'h61EC) & (stage_adr != 2'h3) & ~reg_wait
			 & ~wait_block_brtf ;

// for EVA
        wire            fchram_mask;
        wire            pcwaitf_maccess;
        wire            pcwaitf_pre;
        reg             waitexm_ice;

        // WAITEXM���å��������档PCWAITF����Υޥ����˻��Ѥ��롣
        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb)      waitexm_ice <= 1'b0 ;
                else            waitexm_ice <= waitexm ;
        end

        assign fchram_mask = fchiram & (pc_jump_address[19:16] <= flsize) & (stage_adr == 2'h3) ;

        // �ե��å��Х�����Ѥ���ǡ��������������Ф���PCWAITF��ޥ������롣
        assign pcwaitf_maccess = fchiram_skp | romrd_skp | (slexm & fchiram & dec_ma_enable) ;

        assign pcwaitf_pre = ((pc_wait_flg | pa_st2 | pa_st1 | pa_st0 | waitint) & (stage_adr == 2'h0)) | pcwaitf_maccess |
                             ((stage_adr == 2'h1) & fchiram & pc_wait_flg) | fchram_mask | (fchiram & waitdma) | waitfl ;

        // RAM(EXMEM)�ե��å����EXMEM����������PCWAITF��ޥ������롣�������ե��å����������ϥޥ������ʤ���
        assign pcwaitf = pcwaitf_pre & ~(~fchram & (waitexm | waitexm_ice) & pa_st3) ;

//

// �����������ȿ���Υ������Ȼ��֤򥫥���Ȥ��롣
// ���������ϥ�����ȯ��ľ���RAM�ե��å���Υ�������ȯ��ľ��Υߥ顼�����������ˤϡ�
// �������Ȳ�������ȯ�����ɤ����ᥫ������ͤ��ݻ�����롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)		pc_wait_cnt <= 2'h0 ;
		else if (cpuen) begin
			if (pc_wait_slv)	pc_wait_cnt <= 2'h0 ;
			else if ((data_hazard || (fchiram && (pc_wait_cnt == 2'h1))) && slmirr) pc_wait_cnt <= pc_wait_cnt ;
			else if (pc_wait_flg)	pc_wait_cnt <= pc_wait_cnt + 2'h1 ;
		end
	end

// ������������ȯ��������档���������װ����б���������å����򥫥���Ȥ����飱�ˤʤ롣
	always @(pc_wait_cnt or fchiram_wait or prefix_wait or slmirr) begin
		if (slmirr)		pc_wait_slv = (pc_wait_cnt == 2'h2) ;
		else if (prefix_wait)	pc_wait_slv = (pc_wait_cnt == 2'h2) ;
		else if (fchiram_wait)	pc_wait_slv = (pc_wait_cnt == 2'h2) ;
		else			pc_wait_slv = (pc_wait_cnt == 2'h1) ;
	end

/*------------------------------------------------------------------------------*/
/* �ңϣͥ��ɥ쥹�Υ��󥯥���ȿ��������					*/
/*------------------------------------------------------------------------------*/
/*   �ե��å�������������ңϣͥ��ɥ쥹�Υ��󥯥���Ⱦ���ץ���५����	*/
/*   �β��̣��ӥåȤȸ��߼¹Ԥ��Ƥ���̿���̿��Ĺ���������롣			*/
/*------------------------------------------------------------------------------*/

// PA�Υ��󥯥���Ⱦ�
// PA�򹹿���������������Ƥ��Ƥ⡢�ϥ����ɤ�ȯ�����Ƥ������ϡ�
// PA�ι�����¹Ԥ��ʤ���
	always @(pc or dec_pc_inc1 or dec_pc_inc2 or dec_pc_inc3 or dec_pc_inc4) begin
		casex ({pc[1:0],dec_pc_inc1,dec_pc_inc2,dec_pc_inc3,dec_pc_inc4})
			6'b00_0001 : inc_pa_pre	= 1'b1 ;
			6'b01_0001 : inc_pa_pre	= 1'b1 ;
			6'b01_0010 : inc_pa_pre	= 1'b1 ;
			6'b10_0001 : inc_pa_pre	= 1'b1 ;
			6'b10_0010 : inc_pa_pre	= 1'b1 ;
			6'b10_0100 : inc_pa_pre	= 1'b1 ;
			6'b11_0001 : inc_pa_pre	= 1'b1 ;
			6'b11_0010 : inc_pa_pre	= 1'b1 ;
			6'b11_0100 : inc_pa_pre	= 1'b1 ;
			6'b11_1000 : inc_pa_pre	= 1'b1 ;
			default   : inc_pa_pre = 1'b0 ;
		endcase
	end

	assign	inc_pa = inc_pa_pre & ~data_hazard_flg ;

/*------------------------------------------------------------------------------*/
/* �ңϣͥ��ɥ쥹�Υ��󥯥���Ⱦ���						*/
/*------------------------------------------------------------------------------*/
/*   �ңϣͥ��ɥ쥹�����󥯥���Ȥ��줿�����̿��ʬ�ݻ����롣		*/
/*   �ңϣͥ��ɥ쥹������Ϣ³�ǥ��󥯥���Ȥ��줿���򼨤�������������롣	*/
/*   �����ο���ǡ�̿�ᥭ�塼��ž�����ѥ��ץ饤��ؤ�̿�ᶡ������椹�롣	*/
/*------------------------------------------------------------------------------*/

// ��̿������PA�����󥯥���Ȥ��줿����ɽ�����档
// �ǡ����Х����ɤ������������ȯ�����ȥޥ����������̿��ʳ���FLASH�꡼�ɥ��������ޤ��ϡ�
// RAM�ե��å����FLASH�꡼�ɤȥϥ�����ȯ�������ݻ�����롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)		inc_pa_mst <= 1'b0 ;
		else if (cpuen) begin
			if ((pc_wait_flg && !data_hazard_flg) || (romrd_wait && !(pa_data_mlt1 || pa_data_cyc1)) ||
			   (fchiram && (pa_st2 || data_hazard_flg)))
								inc_pa_mst <= inc_pa_mst ;
			else					inc_pa_mst <= inc_pa ;
		end
	end

// ��̿������PA�����󥯥���Ȥ��줿����ɽ�����档
// ����̿���PA�����󥯥���Ȥ���Ƥ������Υǡ����ϥ����ɤ������������ȯ�����ޤ��ϡ�
// RAM�ե��å����FLASH�꡼�ɤȥϥ�����ȯ�������ݻ�����롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)		inc_pa_slv <= 1'b0 ;
		else if (cpuen) begin
			if ((pc_wait_flg && !(data_hazard_flg && !inc_pa_mst)) || (romrd_wait && !(pa_data_mlt1 || pa_data_cyc1)) ||
			   (fchiram && (pa_st2 | data_hazard_flg)))
								inc_pa_slv <= inc_pa_slv ;
			else					inc_pa_slv <= inc_pa_mst ;
		end
	end

/*------------------------------------------------------------------------------*/
/* �ң��ͥե��å��������������濮��						*/
/*------------------------------------------------------------------------------*/
/*   �ң��ͥե��å���ң��ͥǡ�������������ȯ����̿��ǡ����μ��ľ���򤷤Ƥ���	*/
/*   �֡�̿��μ¹Ԥ򥹥��åפ��롣						*/
/*------------------------------------------------------------------------------*/

// RAM�ե��å����RAM����������ȯ��������磱�Ȥʤ롣
// ̿��¹Ԥ�NOP���֤������륹���å��װ���
	assign fchiram_skp = fchiram & ma_enable_slv ;

/*------------------------------------------------------------------------------*/
/* ̿�������ԥե��å��ѥ��ɥ쥹����						*/
/*------------------------------------------------------------------------------*/
/*   �ץ���५���󥿤��Ф��ƣ�̿��ʬ��Ԥ���̿���ե��å����롣		*/
/*   �ץ���ॢ�ɥ쥹�ȥץ���५���󥿤ε�Υ��׻�����������̿�ᡢ	*/
/*   �ң��ͥե��å���Σң��ͥ����������ңϣͥǡ������������ʤɤǵ�Υ��		*/
/*   �̤ޤä�����ԥե��å���Ԥʤ���						*/
/*   �ץ���ॢ�ɥ쥹�ϥ쥸���������������׼¹Ի��ˤϡ��������襢�ɥ쥹��	*/
/*   ľ�ܽ��Ϥ�ʬ���ڥʥ�ƥ���ڸ����Ƥ��롣					*/
/*------------------------------------------------------------------------------*/

// PA��PC�κ���
	assign	distance_pa_pc = pa_pre[1:0] - pc[3:2] ;

// PA��PC�κ����̾�̿�᤬�¹Ԥ���Ƥ�����Ͼ��3�Ȥʤꡢ�����ס�������ľ��ʤɤ�0����2�Ȥʤ롣
// ��������������̿��¹Ի��������߽����¹Ի���FLASH�꡼�ɥ�����������distance_pa_pc���ͤˤ�餺3�Ȥʤ롣
	assign	pa_inc_en = (pc_jump_en || pa_data_maw || pa_data_buf || pa_data_mlt1 || pa_data_cyc1 || intack_internal) ?
				 2'h3 : distance_pa_pc ;

// PA��PC�ξ��֤�ɽ�����档
	assign	pa_st0 = (pa_inc_en == 2'h0) ;
	assign	pa_st1 = (pa_inc_en == 2'h1) ;
	assign	pa_st2 = (pa_inc_en == 2'h2) ;
	assign	pa_st3 = (pa_inc_en == 2'h3) ;

// ʬ��̿���PC���Ѳ����ᤤ���ᡢ�ץ�ե��å����OCD�μ¹Ը�֥졼����ޥ������롣
	assign	brkmsk = pa_st0 | pa_st1 | pa_st2 ;

// �ץ���ॢ�ɥ쥹���̾��inc_pa�ǥ��󥯥���Ȥ���롣
// FLASH�꡼�ɥ��������ʳ����������������װ����ݻ�����롣
// ������̿��¹Ի��ϡ��������褬RAM���֤��ä����ϥ������襢�ɥ쥹�����Τޤޡ�
// FLASH���֤��ä����ϡ�������å����˥������襢�ɥ쥹�����Ϥ���Ƥ��뤿�ᡢ
// �������襢�ɥ쥹�򥤥󥯥���Ȥ��������ɥ쥹�������ޤ�롣
// RAM�ե��å����RAM��������������դ�������̿�᤬ȯ��������硢PA�ϥǥ�����Ȥ���뤬��
// PA�Υ��󥯥���Ⱦ��ȽŤʤä������ݻ�����롣
// PA���Ե�§�Ѳ����ľ���(pa_jump_en)�Ǥϡ��̾��maw�������ޤ�뤬��
// FLASH�꡼�ɥ���������ȼ��̿�᤬��λ����ݤϡ�RAM�ե��å���Ǥʤ�PA�����󥯥���Ȥ���ʤ���С�
// PC+8����ʳ��ξ��Ǥ�PC+12�������ޤ�롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)
			pa_pre <= 18'h0 ;
		else if (cpuen) begin
			if (!(prefix_wait || slmirr) && pc_wait_flg)
				pa_pre <= pa_pre ;
			else if (pc_jump_en)
				if (((pc_jump_address[19:16] > flsize) & (pc_jump_address[19:10] < {4'hE,2'b11,bfsize})) ||
				     (pc_jump_address[19:16] == 4'hf))
									pa_pre <= pc_jump_address[19:2] ;
				else					pa_pre <= pc_jump_address[19:2] + 18'h00001 ;
			else if (fchiram && !prefix_wait && !slmirr &&
				((dec_ma_enable) && pa_st3 && (dec_clear_stage))) begin
				pa_pre <= pa_pre ;
			end
			else if (pa_jump_en) begin
			// FLASH���ɤߤ�����ˡ�PA���ɤ߽Ф����ξ��֤��᤹��
			// FLASH�꡼�ɥ������󥹤�pa_data_maw�Ǥϡܣ���pa_data_buf�ʹߤǤϡܣ������������ޥ����������̿��Ͻ�����
			// �ޥ����������̿��ξ�硢pa_data_maw�ϡ�High���֤���ӡ��ʹߤο���Ϥ���Ƥ�����
				if ((pa_data_maw || pa_data_buf || pa_data_mlt1 || pa_data_cyc1)) begin
					if (pa_data_maw)	pa_pre <= pc[19:2] + 18'h00002 ;
					else			pa_pre <= pc[19:2] + 18'h00003 ;
				end
				else if (prefix_exe)	pa_pre <= {maw[19:16], maw[15:2]} ;
				else if (slmirr)	pa_pre <= {3'b000, MAA, maw[15:2]} ;
			end
			else if ((pa_inc_en != 2'h3) || inc_pa)
				pa_pre <= pa_pre + 18'h00001 ;
		end
	end

// �ºݤΥץ���ॢ�ɥ쥹��
// ������̿��¹Ի���pc_jump_address��ľ�ܽ��Ϥ���롣
	assign pa = (pc_jump_en) ? pc_jump_address[19:2] : pa_pre ;

// PC��BFLASH��BRAM���֤�ؤ�����磱�Ȥʤ롣
	assign slbmem = ((pc[19:10] >= {4'hE,2'b11,bfsize}) & (pc[19:16] < 4'hF)) ||
			((pc[19:11] >= {4'hF,4'h0,1'b1}) & (pc[19:9] < {4'hF,3'b000,bmsize})) ;

/*------------------------------------------------------------------------------*/
/* �ץ���५����								*/
/*------------------------------------------------------------------------------*/
/*   �ץ���५���󥿤�¹Ԥ��Ƥ���̿���̿��Ĺ�˱����ƥ��󥯥���Ȥ��롣	*/
/*------------------------------------------------------------------------------*/

// �¹Ԥ����̿���̿��Ĺ�˱�����PC�Υ��󥯥�����ͤ�����
	always @(pc or dec_pc_inc1 or dec_pc_inc2 or dec_pc_inc3 or dec_pc_inc4) begin
		if (dec_pc_inc1)	pc_inc = pc + 20'h00001 ;
		else if (dec_pc_inc2)	pc_inc = pc + 20'h00002 ;
		else if (dec_pc_inc3)	pc_inc = pc + 20'h00003 ;
		else if (dec_pc_inc4)	pc_inc = pc + 20'h00004 ;
		else			pc_inc = pc ;
	end

// �ץ���५���󥿡��̾��̿��¹Ծ���(pa_st3)�ǥ��󥯥���Ȥ���롣
// ������̿��¹Ի���pc_jump_address������ࡣ
// FLASH�ե��å����FLASH�꡼�ɼ¹ԤκǸ�ޤ�PC���ݻ����롣
// ��������FLASH�꡼�ɤ��ޥ������������ä����ϡ�slmirr�����Ǥϡ�­��ʤ��Τǡ�pa_data_mlt1��ɬ�ס�
// RAM�ե��å����RAM���������¹ԤκǸ�ޤ�PC���ݻ����롣
// PA�Ȥκ����ͤޤäƤ��ޤ����ץ�ե��å����֤���������ɤ���
// ʬ�����ˤϡ�PC���ݻ����ʤ���
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)						pc <= 20'h0 ;
		else if (cpuen) begin
	 		if (pc_wait_flg || slmirr || prefix_wait || (pa_data_mlt1 & !pc_jump_en) || (fchiram && dec_ma_enable && !pc_jump_en))
									pc <= pc ;
			else if (dec_pc_set_enable && pc_jump_en)	pc <= pc_jump_address ;
			else if (pc_set_op01)				pc <= pc_jump_address ;
			else if (pa_st3)				pc <= pc_inc ;
		end
	end

/*------------------------------------------------------------------------------*/
/* Ver2.0  PC,imdr�Υǡ����饤�󥲡��ƥ��󥰡���ή�︺�Τ����			*/
/*------------------------------------------------------------------------------*/
/* Ver3.0  �ǥ��쥤�ˤ��ҥ��ɻߤ��к���ľ��(CPUV1.5���������᤹)		*/
/*------------------------------------------------------------------------------*/

	assign imdr_groupC = imdr ;
//	assign imdr_groupC = (fchiram) ? imdr : 16'h0000;

/*------------------------------------------------------------------------------*/
/* ̿�ᥭ�塼									*/
/*------------------------------------------------------------------------------*/
/*   ̿����꤫��ե��å�����̿���̿�ᥭ�塼�˽缡ž�����롣			*/
/*------------------------------------------------------------------------------*/
/* Ver2.0��imdr�����Ϥ�imdr_groupC���ѹ�					*/
/*------------------------------------------------------------------------------*/

// RAM�ե��å����̿�ᥭ�塼��ž����郎��Ω������祻�åȤ���롣
// RAM�ե��å���ϡ����塼��ž���ˤ��ο������Ѥ��롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)	inc_que_flg <= 1'b0 ;
		else if (cpuen)	inc_que_flg <= fchiram & (~pa_st3 | inc_pa) ;
	end

// ̿�ᥭ�塼��
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)
			id_que1 <= 32'h0 ;
		else if (cpuen) begin
			if (fchiram) begin
			// RAM�ե��å����̿�ᥭ�塼ž����
			// RAM�Υǡ����˥�����������ݤϡ�̿��ˤ�ä�inc_pa��Ω�äƤ���Τǡ��ݻ���ͥ�褹�롣
				if (ma_enable_fchiram)
					id_que1 <= id_que1 ;
				else if (inc_que_flg) begin
					id_que1[7:0] <= id_que1[23:16] ;
					id_que1[15:8] <= id_que1[31:24] ;
					id_que1[23:16] <= imdr_groupC[7:0] ;
					id_que1[31:24] <= imdr_groupC[15:8] ;
				end
			end
			else begin
			// ROM�ե��å��桢���塼�ϡ�
			// �ޤ��ϥץ�ե��å�����(!pa_st3)���ޤ���PA������(inc_pa)��PID�Υǡ���������ࡣ
			// FLASH�Υǡ������ɤ߽Ф��ݤϡ�̿��ˤ�ä�inc_pa�����ˤʤäƤ���Τǡ��ݻ���ͥ�褹�롣
			// ��������FLASH�꡼�ɤ��ޥ������������ä����ϡ�slmirr�����Ǥϡ�­��ʤ��Τǡ�pa_data_mlt1��ɬ�ס�
			// ʬ�����ˤ��ݻ����ʤ���
				if (slmirr || prefix_wait || (pa_data_mlt1 && !pc_jump_en))
					id_que1 <= id_que1 ;
				else if (!pa_st3 || inc_pa)
					id_que1 <= pid ;
			end
		end
	end

/*------------------------------------------------------------------------------*/
/* �ɣĥ��ơ����Υѥ��ץ饤��쥸����						*/
/*------------------------------------------------------------------------------*/
/*   ̿�ᥭ�塼���ݻ�����Ƥ���̿��ǡ�����ž������̿��Υǥ����ɤ�Ԥʤ���	*/
/*   ���Х��ȤΥ쥸���������Ĥ��ꡢ�¹Ԥ��Ƥ���̿���̿��Ĺ�ˤ��̿�ᥭ�塼��̿	*/
/*   ��ǡ����Х����ޤ��ϴ��˥ѥ��ץ饤��쥸�������ݻ�����Ƥ���ǡ�����ž��	*/
/*   ���롣������̿��¹Ի����ң��ͥե��å���Σң��ͥ�������̿��ľ�塢�ңϣ�	*/
/*   ���������¹Ի��ˤϡ��㳰Ū�˥ǡ����Υ��ꥢ�ޤ����ݻ���Ԥʤ���		*/
/*   �ң��ͥե��å��⡼�ɤǤϡ�̿��ǡ����Х�������˥ǡ����꡼�ɥХ�����	*/
/*   ̿��ǡ�����ž������롣							*/
/*------------------------------------------------------------------------------*/
/* Ver2.0���ǥ�������1stMAP���ˣ��Х����ܤ������ͤ˸��ꤹ�롣			*/
/*�����������ΰ٤�2nd,3rd,4th-MAP���Υǥ����ɿ�������				*/
/*------------------------------------------------------------------------------*/

	assign check234map_10 = (id_que1[7:0] == 8'h31 || id_que1[7:0] == 8'h61 || id_que1[7:0] == 8'h71) ? 1'b1:1'b0;
	assign check234map_11 = (id_que1[15:8] == 8'h31 || id_que1[15:8] == 8'h61 || id_que1[15:8] == 8'h71) ? 1'b1:1'b0;
	assign check234map_12 = (id_que1[23:16] == 8'h31 || id_que1[23:16] == 8'h61 || id_que1[23:16] == 8'h71) ? 1'b1:1'b0;
	assign check234map_13 = (id_que1[31:24] == 8'h31 || id_que1[31:24] == 8'h61 || id_que1[31:24] == 8'h71) ? 1'b1:1'b0;
	assign check234map_01 = (ID_stage1 == 8'h31 || ID_stage1 == 8'h61 || ID_stage1 == 8'h71) ? 1'b1:1'b0;
	assign check234map_02 = (ID_stage2 == 8'h31 || ID_stage2 == 8'h61 || ID_stage2 == 8'h71) ? 1'b1:1'b0;
	assign check234map_03 = (ID_stage3 == 8'h31 || ID_stage3 == 8'h61 || ID_stage3 == 8'h71) ? 1'b1:1'b0;


// for EVA
        assign idpop = dec_sp_inc & ( (ID_stage0[7:4] == 4'hC) | ({ID_stage0,ID_stage1[7:4]} == 12'h61C) ) ;
//

// ID���ơ����Υѥ��ץ饤��쥸�����������˳�Ǽ���줿�ǡ������ǥ����ɤ���롣
// CALLT̿��κݤ˥ơ��֥륢�ɥ쥹������Ǽ���롣�ޤ��������ߤ�̿������ɤ���ʤɤǤϥ��ꥢ����롣
// ������������ȯ������FLASH�꡼�ɥ�����������RAM�ե��å����RAM����������FLASH�꡼�ɥ������������ݻ�����롣
// fchiram_waitȯ�����϶���Ū��MDR�Х��ȣ����ܤΥ��塼����ǡ���������ࡣ
// RAM�ե��å����PREFIX̿��¹Ԥ�RAM���������¹Ը塢̿�����ɤ߾���(pa_st2)��ȯ�����뤬��
// ���ΤȤ���PC���ͤ˱�����MDR�Х���̿�ᥭ�塼����ǡ���������ࡣ
// �ߥ顼���֥�����������PC���ͤ˱����ơ��̾��PID�Х���̿�ᥭ�塼��RAM�ե��å����MDR�Х���̿�ᥭ�塼����ǡ���������ࡣ
// �嵭�ʳ��ξ��ϡ�PC���ͤȼ¹Ԥ����̿���̿��Ĺ�˱����ǥХ��ȣ����ܤΥ��塼�������ܤΥ��塼����ǡ���������ࡣ
// �Х��ϡ��̾�PID�Х�������RAM�ե��å����MDR�Х��Ȥʤ롣
/*------------------------------------------------------------------------------*/
/* Ver2.0���ǥ�������1stMAP���ˣ��Х����ܤ������ͤ˸��ꤹ�롣			*/
/*�����������ΰ٤�ID_stage1_dec�ȥǥ������ѤΣ��Х����ܤΥ쥸��������		*/
/*��������imdr��ɬ�פʻ���������imdr_groupC���ѹ�				*/
/*�����������ɥ쥹���ơ����Υǥ��������Ϥ˥ҥ����Τ뤿�ᡢID_stage0,1����������	*/
/*�������������˥ȥ��뤹��decout_mask_reg����					*/
/*------------------------------------------------------------------------------*/
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) begin
			ID_stage3 <= 8'h00 ;
			ID_stage2 <= 8'h00 ;
			ID_stage1 <= 8'h00 ;
			ID_stage0 <= 8'h00 ;
			ID_stage1_dec <= 8'h00 ;
		end
		else if (cpuen) begin
			if (dec_pc_set_op01) begin
				casex (pc[1])
					1'b1 : ID_stage3 <= pid[31:24] ;
					default : ID_stage3 <= pid[15:8] ;
				endcase
				casex (pc[1])
					1'b1 : ID_stage2 <= pid[23:16] ;
					default : ID_stage2 <= pid[7:0] ;
				endcase
				ID_stage1 <= 8'h00 ;
				ID_stage0 <= 8'h00 ;
				ID_stage1_dec <= 8'h00 ;
			end
			else if (pa_st0 || (pc_set_op01 && !ivack) || pa_st1 || (pc_jump_en && stage_cut_br && !pc_wait_flg) ||
				(dec_pc_set_ret && !pc_wait_flg)) begin
				ID_stage3 <= 8'h00 ;
				ID_stage2 <= 8'h00 ;
				ID_stage1 <= 8'h00 ;
				ID_stage0 <= 8'h00 ;
				ID_stage1_dec <= 8'h00 ;
			end
			// pc_wait_flgȯ�����ˤϡ�ID���ơ����Υ쥸�������ݻ����Ƥ�����
			// FLASH�ե��å����FLASH�꡼�ɻ�(slmirr || prefix_wait)�ˤ��ݻ����롣
			// ��������FLASH�꡼�ɤ��ޥ������������ä����ϡ�slmirr�����Ǥϡ�­��ʤ��Τǡ�pa_data_mlt1��ɬ�ס�
			// RAM�ե��å����RAM����������(fchiram && dec_ma_enable)�ˤ��ݻ����롣
			else if (pc_wait_flg || (pc_jump && !pa_data_cyc1) || ma_enable_fchiram ||
				(!fchiram && (slmirr || prefix_wait || pa_data_mlt1))) begin
				ID_stage3 <= ID_stage3 ;
				ID_stage2 <= ID_stage2 ;
				ID_stage1 <= ID_stage1 ;
				ID_stage0 <= ID_stage0 ;
				ID_stage1_dec <= ID_stage1_dec ;
			end
			else if (fchiram_wait) begin
				ID_stage3 <= imdr_groupC[7:0] ;
				ID_stage2 <= id_que1[31:24] ;
				ID_stage1 <= id_que1[23:16] ;
				ID_stage0 <= id_que1[15:8] ;
				if (check234map_11) ID_stage1_dec <= id_que1[23:16] ;
			end
			else if (fchiram_ramrd || fchiram_romrd) begin
				ID_stage3 <= ID_stage3 ;
				ID_stage2 <= ID_stage2 ;
				ID_stage1 <= ID_stage1 ;
				ID_stage0 <= ID_stage0 ;
				ID_stage1_dec <= ID_stage1_dec ;
			end
			else if (~prefix_ack && pa_st2) begin
				casex ({fchiram,pc[1:0]})
					3'b001 : ID_stage3 <= pid[7:0] ;
					3'b010 : ID_stage3 <= pid[15:8] ;
					3'b011 : ID_stage3 <= pid[23:16] ;
					3'b101 : ID_stage3 <= imdr_groupC[7:0] ;
					3'b110 : ID_stage3 <= imdr_groupC[15:8] ;
					default : ID_stage3 <= id_que1[31:24] ;
				endcase
				casex ({fchiram,pc[1:0]})
					3'bx01 : ID_stage2 <= id_que1[31:24] ;
					3'b010 : ID_stage2 <= pid[7:0] ;
					3'b011 : ID_stage2 <= pid[15:8] ;
					3'b110 : ID_stage2 <= imdr_groupC[7:0] ;
					3'b111 : ID_stage2 <= imdr_groupC[15:8] ;
					default : ID_stage2 <= id_que1[23:16] ;
				endcase
				casex ({fchiram,pc[1:0]})
					3'bx01 : ID_stage1 <= id_que1[23:16] ;
					3'bx10 : ID_stage1 <= id_que1[31:24] ;
					3'b011 : ID_stage1 <= pid[7:0] ;
					3'b111 : ID_stage1 <= imdr_groupC[7:0] ;
					default : ID_stage1 <= id_que1[15:8] ;
				endcase
				casex ({fchiram,pc[1:0]})
					3'bx01 : ID_stage0 <= id_que1[15:8] ;
					3'bx10 : ID_stage0 <= id_que1[23:16] ;
					3'bx11 : ID_stage0 <= id_que1[31:24] ;
					default : ID_stage0 <= id_que1[7:0] ;
				endcase
				casex ({fchiram,pc[1:0]})
					3'bx01 : if (check234map_11) ID_stage1_dec <= id_que1[23:16] ;
					3'bx10 : if (check234map_12) ID_stage1_dec <= id_que1[31:24] ;
					3'b011 : if (check234map_13) ID_stage1_dec <= pid[7:0] ;
					3'b111 : if (check234map_13) ID_stage1_dec <= imdr_groupC[7:0] ;
					default : if (check234map_10) ID_stage1_dec <= id_que1[15:8] ;
				endcase
			end
			else if (dec_pc_inc1) begin
				casex ({fchiram,pc[1:0]})
					3'bx01 : ID_stage3 <= id_que1[15:8] ;
					3'bx10 : ID_stage3 <= id_que1[23:16] ;
					3'bx11 : ID_stage3 <= id_que1[31:24] ;
					default : ID_stage3 <= id_que1[7:0] ;
				endcase
				ID_stage2 <= ID_stage3 ;
				ID_stage1 <= ID_stage2 ;
				ID_stage0 <= ID_stage1 ;
				if (check234map_01) ID_stage1_dec <= ID_stage2;
			end
			else if (dec_pc_inc2) begin
				casex ({fchiram,pc[1:0]})
					3'bx01 : ID_stage3 <= id_que1[23:16] ;
					3'bx10 : ID_stage3 <= id_que1[31:24] ;
					3'b011 : ID_stage3 <= pid[7:0] ;
					3'b111 : ID_stage3 <= imdr_groupC[7:0] ;
					default : ID_stage3 <= id_que1[15:8] ;
				endcase
				casex ({fchiram,pc[1:0]})
					3'bx01 : ID_stage2 <= id_que1[15:8] ;
					3'bx10 : ID_stage2 <= id_que1[23:16] ;
					3'bx11 : ID_stage2 <= id_que1[31:24] ;
					default	: ID_stage2 <= id_que1[7:0] ;
				endcase
				ID_stage1 <= ID_stage3 ;
				ID_stage0 <= ID_stage2 ;
				if (check234map_02) ID_stage1_dec <= ID_stage3;
			end
			else if (dec_pc_inc3) begin
				casex ({fchiram,pc[1:0]})
					3'bx01 : ID_stage3 <= id_que1[31:24] ;
					3'b010 : ID_stage3 <= pid[7:0] ;
					3'b011 : ID_stage3 <= pid[15:8] ;
					3'b110 : ID_stage3 <= imdr_groupC[7:0] ;
					3'b111 : ID_stage3 <= imdr_groupC[15:8] ;
					default : ID_stage3 <= id_que1[23:16] ;
				endcase
				casex ({fchiram,pc[1:0]})
					3'bx01 : ID_stage2 <= id_que1[23:16] ;
					3'bx10 : ID_stage2 <= id_que1[31:24] ;
					3'b011 : ID_stage2 <= pid[7:0] ;
					3'b111 : ID_stage2 <= imdr_groupC[7:0] ;
					default : ID_stage2 <= id_que1[15:8] ;
				endcase
				casex ({fchiram,pc[1:0]})
					3'bx01 : ID_stage1 <= id_que1[15:8] ;
					3'bx10 : ID_stage1 <= id_que1[23:16] ;
					3'bx11 : ID_stage1 <= id_que1[31:24] ;
					default : ID_stage1 <= id_que1[7:0] ;
				endcase
				ID_stage0 <= ID_stage3 ;
				if (check234map_03) begin
					casex ({fchiram,pc[1:0]})
						3'bx01 : ID_stage1_dec <= id_que1[15:8] ;
						3'bx10 : ID_stage1_dec <= id_que1[23:16] ;
						3'bx11 : ID_stage1_dec <= id_que1[31:24] ;
						default : ID_stage1_dec <= id_que1[7:0] ;
					endcase
				end
			end
			else if (dec_pc_inc4) begin
				casex ({fchiram,pc[1:0]})
					3'b001 : ID_stage3 <= pid[7:0] ;
					3'b010 : ID_stage3 <= pid[15:8] ;
					3'b011 : ID_stage3 <= pid[23:16] ;
					3'b101 : ID_stage3 <= imdr_groupC[7:0] ;
					3'b110 : ID_stage3 <= imdr_groupC[15:8] ;
					3'b111 : ID_stage3 <= imdr_groupC[7:0] ;
					default : ID_stage3 <= id_que1[31:24] ;
				endcase
				casex ({fchiram,pc[1:0]})
					3'bx01 : ID_stage2 <= id_que1[31:24] ;
					3'b010 : ID_stage2 <= pid[7:0] ;
					3'b011 : ID_stage2 <= pid[15:8] ;
					3'b110 : ID_stage2 <= imdr_groupC[7:0] ;
					3'b111 : ID_stage2 <= imdr_groupC[15:8] ;
					default : ID_stage2 <= id_que1[23:16] ;
				endcase
				casex ({fchiram,pc[1:0]})
					3'bx01 : ID_stage1 <= id_que1[23:16] ;
					3'bx10 : ID_stage1 <= id_que1[31:24] ;
					3'b011 : ID_stage1 <= pid[7:0] ;
					3'b111 : ID_stage1 <= imdr_groupC[7:0] ;
					default : ID_stage1 <= id_que1[15:8] ;
				endcase
				casex ({fchiram,pc[1:0]})
					3'bx01 : ID_stage0 <= id_que1[15:8] ;
					3'bx10 : ID_stage0 <= id_que1[23:16] ;
					3'bx11 : ID_stage0 <= id_que1[31:24] ;
					default : ID_stage0 <= id_que1[7:0] ;
				endcase
				casex ({fchiram,pc[1:0]})
					3'bx01 : if (check234map_11) ID_stage1_dec <= id_que1[23:16] ;
					3'bx10 : if (check234map_12) ID_stage1_dec <= id_que1[31:24] ;
					3'b011 : if (check234map_13) ID_stage1_dec <= pid[7:0] ;
					3'b111 : if (check234map_13) ID_stage1_dec <= imdr_groupC[7:0] ;
					default : if (check234map_10) ID_stage1_dec <= id_que1[15:8] ;
				endcase
			end
		end
	end

/*------------------------------------------------------------------------------*/
/* �ޥ����������̿�������							*/
/*------------------------------------------------------------------------------*/
/*   �¹Ԥ�ʣ������å���ɬ�פȤ���̿��Υ���å����򼨤���			*/
/*------------------------------------------------------------------------------*/

// ̿��¹��楫����ȥ��åפ��졢��λ����Ω�������롣
// ����ʬ��̿��ϣ�����å��¹ԤʤΤǥ�����ȥ��åפ������Ϥʤ�����
// ������̿���꡼�ɥ�ǥ��ե����饤��̿��Ǥϥ�����ȥ��åפ��롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)					stage_adr <= 2'h0 ;
		else if (cpuen) begin
			if (pc_wait_flg | pa_st2)		stage_adr <= stage_adr ;
			else if (dec_clear_stage | brunch_en)	stage_adr <= 2'h0 ;
			else					stage_adr <= stage_adr + 2'h1 ;
		end
	end

/*------------------------------------------------------------------------------*/
/* �ͣţͥ��ơ����Υѥ��ץ饤��쥸����						*/
/*------------------------------------------------------------------------------*/
/*   �ɣĥ��ơ������饪�ڥ��ɥǡ�����ž������롣���Х��ȤΥ쥸�������Ĥ�	*/
/*   �������졢���̣դˤ��黻��ɬ�פʥ��ڥ��ɤΤߤ�ž������롣		*/
/*------------------------------------------------------------------------------*/

// MEM���ơ����Υѥ��ץ饤��쥸���������Υǡ��������ڥ��ɤȤ��Ʊ黻�ʤɤ˻��Ѥ���롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) begin
			MEM_stage0 <= 8'h00 ;
		end
		else if (cpuen) begin
			if (dec_mem_stage_op2)		MEM_stage0 <= ID_stage2 ;
			else if (dec_mem_stage_op3)	MEM_stage0 <= ID_stage3 ;
			else if (dec_mem_stage_op23)	MEM_stage0 <= ID_stage2 ;
			else				MEM_stage0 <= ID_stage1 ;
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) begin
			MEM_stage1 <= 8'h00 ;
		end
		else if (cpuen) begin
			if (dec_mem_stage_op23)		MEM_stage1 <= ID_stage3 ;
			else				MEM_stage1 <= ID_stage2 ;
		end
	end

/*------------------------------------------------------------------------------*/
/* �ǡ����ϥ����ɥե饰								*/
/*------------------------------------------------------------------------------*/
/*   ���ѥ쥸�����ؤΥ����������ɣĥ��ơ����ȣͣţͥ��ơ����ǽ�ʣ������硢	*/
/*   �ǡ����ϥ����ɥե饰���������롣						*/
/*   �ң��ͥե��å��������������ңϣͥǡ������������������ѥ쥸�����ؤ�������	*/
/*   �ǡ���ž����ޥ������롣���������ң��ͥե��å���˥ϥ�����ȯ����������	*/
/*   ��������ư���ͭ���뤿�ᡢ�㳰Ū��ž������Ĥ��롣			*/
/*------------------------------------------------------------------------------*/

// �쥸�����ڥ������򤵤줿��磱�Ȥʤ롣
	assign pc_set_rp = dec_pc_set_AX | dec_pc_set_BC | dec_pc_set_DE | dec_pc_set_HL ;

// SP�����ȳ����ߤ�ޤ�ʬ��̿��Ȥ�Hazardȯ�����ˣ��Ȥʤ롣
// RAM�ե��å��¹�����ü�����椬ɬ�פʤ��ᡢ¾�Υϥ������װ��ȶ��̤��롣
	assign sp_hazard_flg = (dec_ma_data_sp | dec_ma_data_SPop1 | dec_sp_set_enable) & SP_enable ;

// �ǡ����ϥ�����ȯ���ե饰��
// ���ѥ쥸�����ؤν񤭹���̿���MEM���ơ����ȥ쥸�������ɥ�å��󥰤ޤ��ϥ����å�ư���ID���ơ�����
// Ʊ���쥸�����Ǥ֤Ĥ��ä���磱�Ȥʤ롣
// �ޤ��Х��ڤ��ؤ�̿�ᡢPSW���������ȥ쥸�����ˤ����ܥ��ꥢ���������֤Ĥ��ä����⣱�Ȥʤ롣
	assign data_hazard_flg_pre = ((dec_ma_data_DE | dec_ma_data_DEop1 | dec_ma_data_DEop2)
										&	(D_access | E_access | dec_RBS_enable)) |
				     ((dec_ma_data_HL | dec_ma_data_HLop1 | dec_ma_data_HLop2 | dec_ma_data_HLB | dec_ma_data_HLC)
										&	(H_access | L_access | dec_RBS_enable)) |
				      (dec_ma_data_BCop12			&	(B_access | C_access | dec_RBS_enable)) |
				     ((dec_ma_data_Bop12 | dec_ma_data_HLB)	&	(B_access | dec_RBS_enable)) |
				     ((dec_ma_data_Cop12 | dec_ma_data_HLC)	&	(C_access | dec_RBS_enable)) |
				      sp_hazard_flg |
				     (dec_pc_set_AX				&	(A_access | X_access | dec_RBS_enable)) |
				     (dec_pc_set_BC				&	(B_access | C_access | dec_RBS_enable)) |
				     (dec_pc_set_DE				&	(D_access | E_access | dec_RBS_enable)) |
				     (dec_pc_set_HL				&	(H_access | L_access | dec_RBS_enable)) |
				     (pc_set_rp					&	CS_enable) ;

// RAM�ե��å��ˤ�륦��������ϡ��ϥ����ɾ�郎��Ω���Ƥ�̵���Ȥ��롣
	assign data_hazard_flg = data_hazard_flg_pre & ~(fchiram & (pc_wait_cnt != 0)) ;

// ������å����˥ϥ����ɤ�ȯ����������ɽ�����档
// RAM�ե��å����Ω���ʤ���
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) data_hazard <= 1'b0 ;
		else if (cpuen) begin
			if (fchiram) data_hazard <= 1'b0 ;
			else data_hazard <= data_hazard_flg ;
		end
	end

// ������å�����SP�ˤ��ϥ����ɤ�ȯ����������ɽ������
// RAM�ե��å���Τߣ��ȤʤꡢMA��SP�ι�������Ĥ��롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) sp_hazard <= 1'b0 ;
		else if (cpuen) begin
			if (sp_hazard) sp_hazard <= 1'b0 ;
			else sp_hazard <= sp_hazard_flg & fchiram ;
		end
	end

// RAM�ե��å����Flash�꡼�ɥ���������ˡ��쥸�����Υǡ������ݻ����뤿��ο��档
	assign reg_wait = ~(data_hazard_flg) &
			 ((fchiram & (pc_wait_cnt != 0)) |
			 pa_data_maw | pa_data_buf )  ;

/*------------------------------------------------------------------------------*/
/* �ꥻ�åȥ٥����ե饰								*/
/*------------------------------------------------------------------------------*/
/*   �ꥻ�åȥ٥����ե饰���������롣						*/
/*------------------------------------------------------------------------------*/

// PC�����Ǥ��ä���磱�Ȥʤ롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) rstvec <= 1'b0 ;
		else if (cpuen) begin
			if (rstvec || pc_set_op01) rstvec <= 1'b0 ;
// for EVA
//			else if (pc == 20'h0) rstvec <= 1'b1 ;
                        else if ((pc == 20'h0) & !svmod) rstvec <= 1'b1 ;
//
		end
	end

/*------------------------------------------------------------------------------*/
/* �����߼����դ��ե饰							*/
/*------------------------------------------------------------------------------*/
/*   ̿��¹���ޤ��ϡ���������α̿���ɣťե饰��Ƚ�̤��������߼����դ�	*/
/*   �ե饰���������롣								*/
/*------------------------------------------------------------------------------*/

// �ޥ����֥�����߼¹Զػ߿��档PSW��������磱�Ȥʤꡢ�����߼¹Ԥ϶ػߤȤʤ롣
// DMAž�������դ����ˤ⣱�Ȥ������inten��Ω�������롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)				inten_block <= 1'b0 ;
		else if (cpuen) begin
			if (pc_wait_flg && !fchiram)	inten_block <= inten_block ;
			else if ((reg_wait || (pa_st2 && pc_wait_flg)) && fchiram)	inten_block <= inten_block ;
			else if (pa_st3 || pa_st2)	inten_block <= PSW_block & dec_cpuwr_enable ;
		end
	end

// �Υ�ޥ����֥�����߼¹Զػ߿��档PSW��������磱�Ȥʤꡢ�����߼¹Ԥ϶ػߤȤʤ롣
// DMAž�������դ����ˤ⣱�Ȥ������inten��Ω�������롣RAM�ե��å����High���ֱ�Ĺ��
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) 				nmien_block <= 1'b0 ;
		else if (cpuen) begin
			if (pc_wait_flg && !fchiram)	nmien_block <= nmien_block ;
			else if ((reg_wait || (pa_st2 && pc_wait_flg)) && fchiram)	nmien_block <= nmien_block ;
			else if (pa_st3 || pa_st2)	nmien_block <= (dec_pc_set_ret & intblock) | dmaack ;
		end
	end

// �ޥ����֥��������α���档
// PSW��������硢INT�ޥ����SFR��������硢PUSH/POP PSW̿��ϳ������׵᤬��α����롣
// DMA�����դ����ˤ�����ߤ���α����롣DMA�׵�ȳ������׵᤬Ʊ���Ǥ����DMA��ͥ�褵��롣
// ��������RAM�ե��å����RAM��������ľ��˸¤äƤϡ�ID���ơ����Ǥγ�������α��̵�������롣
	assign int_suspend = inten_block | nmien_block |
			(
			( ( (PSW_block | (maw == 20'hffffa) | ((maw[19:4] == 16'hfffe) | (maw[19:4] == 16'hfffd))) & dec_cpuwr_enable ) |
			({ID_stage0,ID_stage1} == 16'h61CD)) & ~(fchiram_skp | romrd_skp)
			) ;

// RAM�ե��å���Υ��ꥢ������ư�λ�ޤǳ�������α������ݻ����Ƥ�����
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) 			int_suspend_fchiram <= 1'b0 ;
		else if (cpuen) begin
			if (pc_wait_flg)	int_suspend_fchiram <= int_suspend_fchiram ;
			else			int_suspend_fchiram <= int_suspend & fchiram & dec_ma_enable;
		end
	end

// �Υ�ޥ����֥��������α���档
// DMA�����դ����ˤ�����ߤ���α����롣DMA�׵�ȳ������׵᤬Ʊ���Ǥ����DMA��ͥ�褵��롣
// for EVA
//	assign nmi_suspend = nmien_block | ((ID_stage0 == 8'h11) & ~(fchiram_skp | romrd_skp)) |
//			     skp_block | dmaack | (dmarq & ~(intdbg | intnmi)) ;
        assign nmi_suspend = svmod | nmien_block | ((ID_stage0 == 8'h11) & ~(fchiram_skp | romrd_skp)) |
                             skp_block | dmaack | (dmarq & ~(intdbg | intnmi | svi)) ;
//

// �����߼����դ���ǽ���֤ǣ��Ȥʤ롣
// ��������α̿��Ǥʤ���̿��¹�����Ǥʤ���г����߼����դ���ǽ��
// �ޥ����֥롿�Υ�ޥ����֥���鷺���ο��椬���Ǥʤ���г����ߤϼ����դ��ʤ���
	assign iopen = (pa_st3 | pa_st2) & (dec_clear_stage | pa_data_mem) & ~pc_wait_flg & ~(fchiram & dec_ma_enable) &
			~(pc_jump_en | pa_data_maw | pa_data_buf | pa_data_mlt1 | pa_data_cyc1 | intack_internal) ;

// �����ߵ��ľ��֤Ǥ��ĥޥ����֥�����߼����դ���ǽ�Ǥ���У��Ȥʤ롣
	assign inten = IE & iopen & ~int_suspend & ~nmi_suspend & ~int_suspend_fchiram ;

// �Υ�ޥ����֥�����߼����դ���ǽ�Ǥ���У��Ȥʤ롣
	assign nmien = iopen & ~nmi_suspend ;

/*------------------------------------------------------------------------------*/
/* ������ͥ����Ƚ��								*/
/*------------------------------------------------------------------------------*/
/*   �ޥ����֥�����ߤ�ͥ���̤�Ƚ�ꤷ�ɣӣХե饰���������롣		*/
/*   �Υ�ޥ����֥롢�ǥХå������ߤ�ͥ���̤�Ƚ�ꤷ���Σͣɣӡ��ģ£ǣ�	*/
/*   �ե饰���������롣								*/
/*   �����߲�ǽ�Ǥ���С�������ư��򳫻Ϥ��롣				*/
/*------------------------------------------------------------------------------*/

/*------------------------------------------------------------------------------*/
/* Ver2.0  ��ή�︺�ΰ١�������׵�ʤ��λ��˳����������ϩ����ߤ��롣	*/
/*------------------------------------------------------------------------------*/
	assign intclk_on = intdbg | intnmi | (IE & (intrq3 | intrq2 | intrq1 | intrq0))  |
			   ivack | dec_NMIS_enable | dec_pc_set_dbg | monmd |
			   svi | svintack | svmod | svmodi | alt1 | alt2;

// �������׵΅��˱�����ISP�ե饰�˼�����٤��ǡ��������򤹤롣
	always @(intrq3 or intrq2 or intrq1 or intrq0) begin
		casex ({intrq3,intrq2,intrq1,intrq0})
			4'b1000 : intisp_pre = 2'b10 ;
			4'b0100 : intisp_pre = 2'b01 ;
			4'b0010 : intisp_pre = 2'b00 ;
			default : intisp_pre = 2'b00 ;
		endcase
	end

// �������׵᤬�����դ���줿��硢���Υǡ�����ISP�ե饰�˳�Ǽ����롣
/*------------------------------------------------------------------------------*/
/* Ver2.0  intclk_on�ǥ����ƥ���						*/
/*------------------------------------------------------------------------------*/
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) intisp <= 2'b00 ;
		else if (cpuen & intclk_on) begin
			if (data_hazard)	intisp <= intisp ;
			else			intisp <= intisp_pre ;
		end
	end

// ͥ���̤�Ƚ�̤����ޥ����֥�����߼����դ���ǽ�ʾ�磱�Ȥʤ롣
/*------------------------------------------------------------------------------*/
/* Ver2.0  intclk_on�ǽ����Ѳ�							*/
/*------------------------------------------------------------------------------*/
	always @(intrq3 or intrq2 or intrq1 or intrq0 or isp or inten or DBGS or NMIS or intclk_on) begin
		if (inten & intclk_on) begin
			casex ({intrq3,intrq2,intrq1,intrq0,isp,DBGS,NMIS})
				8'b1000_11_00 : mkiack = 1'b1 ;
				8'b0100_1x_00 : mkiack = 1'b1 ;
				8'b0010_1x_00 : mkiack = 1'b1 ;
				8'b0010_01_00 : mkiack = 1'b1 ;
				8'b0001_xx_00 : mkiack = 1'b1 ;
				default : mkiack = 1'b0 ;
			endcase
		end
		else	mkiack = 1'b0 ;
	end

// ͥ���̤�Ƚ�ꤷ���Υ�ޥ����֥�����߼����դ���ǽ�ʾ�磱�Ȥʤ롣
// �ޤ����ǥХå������ߥե饰�ȥΥ�ޥ����֥�����ߥե饰�Υǡ��������򤹤롣
// for EVA
//	always @(intdbg or intnmi or DBGS or NMIS or nmien) begin
//		if (nmien) begin
//			casex ({intdbg,intnmi,DBGS,NMIS})
//				4'b1x_0x : {nmiack,dbgd,nmid} = 3'b1_10 ;
//				4'b01_00 : {nmiack,dbgd,nmid} = 3'b1_01 ;
//				default : {nmiack,dbgd,nmid} = 3'b0_00 ;
//			endcase
//		end
//		else	{nmiack,dbgd,nmid} = 3'b0_00 ;
//	end

        wire intnmi_eva = intnmi & ~icemsknmi ;
        wire intdbg_eva = intdbg & ~icemskdbg ;

            always @(intdbg_eva or intnmi_eva or DBGS or NMIS or nmien) begin
                    if (nmien) begin
                            casex ({intdbg_eva,intnmi_eva,DBGS,NMIS})
                                    4'b1x_0x : {nmiack,dbgd,nmid} = 3'b1_10 ;
                                    4'b01_00 : {nmiack,dbgd,nmid} = 3'b1_01 ;
                                    default : {nmiack,dbgd,nmid} = 3'b0_00 ;
                            endcase
                    end
                    else        {nmiack,dbgd,nmid} = 3'b0_00 ;
            end
//
// for EVA

        always @(svi or nmien) begin
                if (nmien) begin
                        sviack = svi ;
                end
                else    sviack = 1'b0 ;
        end

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb)              svintack <= 1'b0 ;
                else if (cpuen) begin
                        if (svintack)   svintack <= 1'b0 ;
                        else            svintack <= sviack ;
                end
        end

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb) begin
                        sviack_buf <= 1'b0 ;
                end
                else if (cpuen) begin
                        if (pc_wait_flg) begin
                                sviack_buf <= sviack_buf ;
                        end
                        else begin
                                sviack_buf <= sviack ;
                        end
                end
        end
//

// �����߼����դ�����򣱥���å��ݻ���ivack��HIGH�����Ĺ���롣
/*------------------------------------------------------------------------------*/
/* Ver2.0  intclk_on�ǥ����ƥ���						*/
/*------------------------------------------------------------------------------*/
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) begin
			nmiack_buf <= 1'b0 ;
			mkiack_buf <= 1'b0 ;
		end
		else if (cpuen & intclk_on) begin
			if (pc_wait_flg) begin
				nmiack_buf <= nmiack_buf ;
				mkiack_buf <= mkiack_buf ;
			end
			else begin
				nmiack_buf <= nmiack ;
				mkiack_buf <= mkiack ;
			end
		end
	end

// �ǥХå������ߡ��Υ�ޥ����֥�����ߥե饰��
// �Υ�ޥ����֥�����߼����դ��塢�ǡ����������ޤ�롣
// �̾�NMIS��RET̿��ǥ��ꥢ����뤬���ǥХå���������ϥ��ꥢ����ʤ���
/*------------------------------------------------------------------------------*/
/* Ver2.0  intclk_on�ǥ����ƥ���						*/
/*------------------------------------------------------------------------------*/
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) begin
			DBGS <= 1'b0 ;
			NMIS <= 1'b0 ;
		end
		else if (cpuen & intclk_on) begin
			if (dec_pc_set_dbg) begin
				DBGS <= 1'b1 ;
			end
			else if (nmiack) begin
				DBGS <= dbgd ;
				NMIS <= nmid ;
			end
			else if (dec_NMIS_enable) begin
				if (!DBGS) begin
					DBGS <= DBGS ;
					NMIS <= 1'b0 ;
				end
				else begin
					DBGS <= 1'b0 ;
					NMIS <= NMIS ;
				end
			end
		end
	end

// �����߱������档�����ߤ������դ���줿��磱�Ȥʤ롣
// �������������߶��祦�����ȡ��������ꥢ����������������ϣ��Ȥ��롣
/*------------------------------------------------------------------------------*/
/* Ver2.0  intclk_on�ǥ����ƥ���						*/
/*------------------------------------------------------------------------------*/
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)		intack_pre <= 1'b0 ;
		else if (cpuen & intclk_on) begin
			if (intack_internal)	intack_pre <= 1'b0 ;
			else		intack_pre <= mkiack | nmiack ;
		end
	end

// for EVA
//
//	assign intack = intack_pre & ~waitint & ~waitexm & ~wait2ndsfr & ~waitfl & ~waitmod ;
//	assign intack = intack_pre & ~waitint & ~waitexm & ~wait2ndsfr & ~waitfl & ~waitmod & ~svintack ;
	assign intack_internal = intack_pre & ~waitint & ~waitexm & ~wait2ndsfr & ~waitdflash & ~waitfl & ~waitmod & ~svintack ;
//	assign intack = intack_internal & ~(RVEON & ~wed) ;
	assign intack = intack_internal & (~(RVEON & ~wed) | (intdbg | dec_pc_set_dbg | hazard_dbgintack)) ;
//

// intack�������ivack��HIGH�����Ĺ���롣
/*------------------------------------------------------------------------------*/
/* Ver2.0  intclk_on�ǥ����ƥ���						*/
/*------------------------------------------------------------------------------*/
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)		ivack_pre <= 1'b0 ;
		else if (cpuen & intclk_on) begin
			if (ivack_pre)	ivack_pre <= 1'b0 ;
// for EVA
//			else		ivack_pre <= intack_internal ;
                        else            ivack_pre <= intack_internal | svintack ;
//
		end
	end

// ivack_pre�������ivack��HIGH�����Ĺ���롣
/*------------------------------------------------------------------------------*/
/* Ver2.0  intclk_on�ǥ����ƥ���						*/
/*------------------------------------------------------------------------------*/
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)		ivack_end <= 1'b0 ;
		else if (cpuen & intclk_on) begin
			if (ivack_end)	ivack_end <= 1'b0 ;
			else		ivack_end <= ivack_pre ;
		end
	end

// �����߽����¹ԥե饰���ǥ������Ϥ��ο���ǳ����߽��������濮����������롣
/*------------------------------------------------------------------------------*/
/* Ver2.0  intclk_on�ǥ����ƥ���						*/
/*------------------------------------------------------------------------------*/
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)		ivack <= 1'b0 ;
// for EVA
//		else if (cpuen & intclk_on)	ivack <= mkiack | nmiack | ivack_pre | ivack_end | nmiack_buf | mkiack_buf ;
                else if (cpuen & intclk_on)     ivack <= sviack | sviack_buf | mkiack | nmiack | ivack_pre | ivack_end | nmiack_buf | mkiack_buf ;
//
	end

// �ϥ�����ȯ�����ˡ��ǥХå������ߤ�INTACK���ݻ����Ƥ�����
/*------------------------------------------------------------------------------*/
/* Ver2.0  intclk_on�ǥ����ƥ���						*/
/*------------------------------------------------------------------------------*/
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)		hazard_dbgintack <= 1'b0 ;
		else if (cpuen & intclk_on) begin
					hazard_dbgintack <= intack_internal & intdbg & data_hazard_flg ;
		end
	end

// for EVA

        // �ϥ�����ȯ������SVINTACK���ݻ����Ƥ���
        reg             hazard_svintack;

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb)              hazard_svintack <= 1'b0 ;
                else if (cpuen) begin
                                        hazard_svintack <= svintack & data_hazard_flg ;
                end
        end
//

// �ǥХå������ߤ������դ���줿����SOFTBREAK���¹Ԥ��줿����Ω���夬�ꡣ
// RETI�ޤ���RETB��Ω�������롣������RETB�ˤ�륯�ꥢ�϶ػߤ����٤���
/*------------------------------------------------------------------------------*/
/* Ver2.0  intclk_on�ǥ����ƥ���						*/
/*------------------------------------------------------------------------------*/
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)					monmd_pre <= 1'b0 ;
		else if (cpuen & intclk_on) begin
// for EVA Ver1.51 OCDMOD�ǡ�OCD�֥졼���桢SVMOD����RETI�����Ȥ���MONMOD����Ȥ��ʤ��褦�ˤ��롣
//			if (pa_st2 && nmien_block && !(fchiram && pc_wait_flg))		monmd_pre <= 1'b0 ;
                        if ((pa_st2 && nmien_block && !(fchiram && pc_wait_flg) && !(ocdmod && svmod))) monmd_pre <= 1'b0 ;
//
			else if (!monmd && data_hazard_flg)	monmd_pre <= 1'b0 ;
// for Eva Ver1.52 monmd��ICE��SoftBreak�Ǥ�Ω�Ƥʤ�
//			else if (monmd || dec_pc_set_dbg)	monmd_pre <= 1'b1 ;
                        else if ((monmd || dec_pc_set_dbg) && ocdmod)   monmd_pre <= 1'b1 ;
// for Eva Ver1.52 modmd��ICE��HardBreak�Ǥ�Ω�Ƥʤ�
			else					monmd_pre <= (intack_internal & intdbg) | hazard_dbgintack ;
		end
	end

// ��˥��⡼�ɿ��档
	assign monmd = monmd_pre ;

// �ǥХå������ߤ������դ���줿����SOFTBREAK���¹Ԥ��줿����Ω���夬�ꡣ
// RETI��Ω�������롣
/*------------------------------------------------------------------------------*/
/* Ver2.0  intclk_on�ǥ����ƥ���						*/
/*------------------------------------------------------------------------------*/
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)					monmdstp_pre <= 1'b0 ;
		else if (cpuen & intclk_on) begin
			// MONMDSTP��RETI�ǤΤ�Ω��������
// for EVA Ver1.51 OCDMOD�ǡ�OCD�֥졼���桢SVMODF����RETI�����Ȥ���MONMODSTP����Ȥ��ʤ��褦�ˤ��롣
//			if (dec_NMIS_enable)			monmdstp_pre <= 1'b0 ;
                        if (dec_NMIS_enable && !(ocdmod && svmodf))     monmdstp_pre <= 1'b0 ;
//
			else if (!monmdstp && data_hazard_flg)	monmdstp_pre <= 1'b0 ;
// for Eva Ver1.52 monmdstp��ICE��SoftBreak�Ǥ�Ω�Ƥʤ�
//			else if (monmdstp || dec_pc_set_dbg)	monmdstp_pre <= 1'b1 ;
                        else if ((monmdstp || dec_pc_set_dbg) && ocdmod)        monmdstp_pre <= 1'b1 ;
// for Eva Ver1.52 modmd��ICE��HardBreak�Ǥ�Ω�Ƥʤ�
			else					monmdstp_pre <= (intack_internal & intdbg) | hazard_dbgintack ;
//
		end
	end

// OCD���ƥå׼¹��ѥ�˥����⡼�ɿ��档
	assign monmdstp = monmdstp_pre ;

// for EVA

        reg             svmod_pre, svmodf_pre, svmodi_pre;

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb)                                      svmod_pre <= 1'b0 ;
                else if (cpuen) begin
                        if (pa_st2 && nmien_block && !(fchiram && pc_wait_flg))         svmod_pre <= 1'b0 ;
                        else if (!svmod && data_hazard_flg)     svmod_pre <= 1'b0 ;
                        else if (svmod)                         svmod_pre <= 1'b1 ;
                        else if (svmod_pre)                     svmod_pre <= 1'b1 ;
                        // Ver1.51
                        //else if (dec_pc_set_dbg)              svmod_pre <= 1'b1 ;
                        else if (dec_pc_set_dbg && !ocdmod)     svmod_pre <= 1'b1 ;
                        else                                    svmod_pre <= svintack | hazard_svintack ;
                end
        end

        assign svmod = svmod_pre ;

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb)                              svmodf_pre <= 1'b0 ;
                else if (cpuen) begin
                        if (!svmodf && data_hazard_flg) svmodf_pre <= 1'b0 ;
                        // Ver1.51
                        //else if (svintack || hazard_svintack || dec_pc_set_dbg)       svmodf_pre <= 1'b1 ;
                        else if (svintack || hazard_svintack || (dec_pc_set_dbg && !ocdmod))    svmodf_pre <= 1'b1 ;
                        // SVMODF��RETI�ǤΤ�Ω��������
                        else if (dec_NMIS_enable)       svmodf_pre <= 1'b0 ;
                        else                            svmodf_pre <= svmodf ;
                end
        end

        // SVMODF�����եȥ֥졼�����ˣ�����å��᤯Ω���夬�롣
        // Ver1.51
        //assign svmodf = svmodf_pre | (dec_pc_set_dbg & ~data_hazard_flg) ;
        assign svmodf = svmodf_pre | ((dec_pc_set_dbg & !ocdmod) & ~data_hazard_flg) ;

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb)              svmodi_pre <= 1'b0 ;
                else if (cpuen) begin
                        if (data_hazard_flg)    svmodi_pre <= svmodi_pre ;
                        else                    svmodi_pre <= sviack ;
                end
        end

        // SP�ȥ����SVMOD���⣱����å��᤯SV�꥽�������ڤ��ؤ���
        // Ver1.51
        //assign svmodi = (svmodi_pre | dec_pc_set_dbg) & ~data_hazard_flg ;
        assign svmodi = (svmodi_pre | (dec_pc_set_dbg & !ocdmod)) & ~data_hazard_flg ;
//

// SOFTBREAK�ǥ�˥��⡼�ɤ����ä����򼨤�������å����ο��档
// �ǥХå������ߤˤ��֥졼���ȶ��̤��뤿����Ѥ��롣
// �ϥ�����ȯ�����ϣ�����å��٤��Ω���夬�롣
/*------------------------------------------------------------------------------*/
/* Ver2.0  intclk_on�ǥ����ƥ���						*/
/*------------------------------------------------------------------------------*/
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)				softbrk <= 1'b0 ;
		else if (cpuen & intclk_on) begin
			if (softbrk)			softbrk <= 1'b0 ;
			else				softbrk <= dec_pc_set_dbg & ~data_hazard_flg ;
		end
	end

/*------------------------------------------------------------------------------*/
/* �ģͣ������դ��ե饰								*/
/*------------------------------------------------------------------------------*/
/*   �ģͣ��׵΅���Ƚ�ꤷ���ģͣ������դ��ե饰���������롣			*/
/*------------------------------------------------------------------------------*/

// PREFIX̿��¹Ի��ˣ��Ȥʤ�DMA���դ���α���롣
	assign dma_suspend = (ID_stage0 == 8'h11) & ~(fchiram_skp | romrd_skp) ;

// DMA�����դ���ǽ���֤ǣ��Ȥʤ롣
// HALT̿��ʳ���̿��¹�����Ǥʤ����DMA�����դ���ǽ��
	assign dopen = ((pa_st3 | pa_st2) & (dec_clear_stage | hltst) & ~pc_wait_flg &
			~(pc_jump_en | pa_data_maw | pa_data_buf | pa_data_mlt1 | pa_data_cyc1 | intack_internal)) & ~dma_suspend ;

// for EVA

        reg             alt1, alt2_pre, alt2;

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb)              alt1i <= 1'b0 ;
                else if (cpuen) begin
                        if (pa_st2)     alt1i <= 1'b0 ;
                        else            alt1i <= dec_alt1 ;
                end
        end

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb)                                      alt1 <= 1'b0 ;
                else if (cpuen) begin
                        if (pa_st2)                             alt1 <= alt1i ;
                        else if (stage_adr != 2'b00)            alt1 <= alt1 ;
                        else if (pa_data_pre)                   alt1 <= alt1 ;
                        else                                    alt1 <= alt1i ;
                end
        end

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb)              alt2_pre <= 1'b0 ;
                else if (cpuen) begin
                                        alt2_pre <= dec_alt2 ;
                end
        end

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb)              alt2 <= 1'b0 ;
                else if (cpuen) begin
                                        alt2 <= alt2_pre ;
                end
        end
//

/*------------------------------------------------------------------------------*/
/* Ver3.0  ���ɥ쥹�Х��Υ����ƥ��󥰲�ϩ�ɲ�					*/
/*         MF2�ޤǤ�OCD�ޥ���Ǽ»ܤ��Ƥ������������ƥ��󥰸�Υ��ɥ쥹��	*/
/*         ���Ѥ���ޥ���򿷵��ɲäΤ���CPU��ǰ�礷�Ƽ»ܤ��롣		*/
/*------------------------------------------------------------------------------*/

	assign	gatead = gatead1 | gatead2 | gatead3 ;

	assign	monpc[19] = gatead & pc[19];
	assign	monpc[18] = gatead & pc[18];
	assign	monpc[17] = gatead & pc[17];
	assign	monpc[16] = gatead & pc[16];
	assign	monpc[15] = gatead & pc[15];
	assign	monpc[14] = gatead & pc[14];
	assign	monpc[13] = gatead & pc[13];
	assign	monpc[12] = gatead & pc[12];
	assign	monpc[11] = gatead & pc[11];
	assign	monpc[10] = gatead & pc[10];
	assign	monpc[9] = gatead & pc[9];
	assign	monpc[8] = gatead & pc[8];
	assign	monpc[7] = gatead & pc[7];
	assign	monpc[6] = gatead & pc[6];
	assign	monpc[5] = gatead & pc[5];
	assign	monpc[4] = gatead & pc[4];
	assign	monpc[3] = gatead & pc[3];
	assign	monpc[2] = gatead & pc[2];
	assign	monpc[1] = gatead & pc[1];
	assign	monpc[0] = gatead & pc[0];

	assign	monma[15] = gatead & ma[15];
	assign	monma[14] = gatead & ma[14];
	assign	monma[13] = gatead & ma[13];
	assign	monma[12] = gatead & ma[12];
	assign	monma[11] = gatead & ma[11];
	assign	monma[10] = gatead & ma[10];
	assign	monma[9] = gatead & ma[9];
	assign	monma[8] = gatead & ma[8];
	assign	monma[7] = gatead & ma[7];
	assign	monma[6] = gatead & ma[6];
	assign	monma[5] = gatead & ma[5];
	assign	monma[4] = gatead & ma[4];
	assign	monma[3] = gatead & ma[3];
	assign	monma[2] = gatead & ma[2];
	assign	monma[1] = gatead & ma[1];
	assign	monma[0] = gatead & ma[0];

	assign	monmdr[15] = gatead & imdr[15];
	assign	monmdr[14] = gatead & imdr[14];
	assign	monmdr[13] = gatead & imdr[13];
	assign	monmdr[12] = gatead & imdr[12];
	assign	monmdr[11] = gatead & imdr[11];
	assign	monmdr[10] = gatead & imdr[10];
	assign	monmdr[9] = gatead & imdr[9];
	assign	monmdr[8] = gatead & imdr[8];
	assign	monmdr[7] = gatead & imdr[7];
	assign	monmdr[6] = gatead & imdr[6];
	assign	monmdr[5] = gatead & imdr[5];
	assign	monmdr[4] = gatead & imdr[4];
	assign	monmdr[3] = gatead & imdr[3];
	assign	monmdr[2] = gatead & imdr[2];
	assign	monmdr[1] = gatead & imdr[1];
	assign	monmdr[0] = gatead & imdr[0];

	assign	monmdw[15] = gatead & mdw[15];
	assign	monmdw[14] = gatead & mdw[14];
	assign	monmdw[13] = gatead & mdw[13];
	assign	monmdw[12] = gatead & mdw[12];
	assign	monmdw[11] = gatead & mdw[11];
	assign	monmdw[10] = gatead & mdw[10];
	assign	monmdw[9] = gatead & mdw[9];
	assign	monmdw[8] = gatead & mdw[8];
	assign	monmdw[7] = gatead & mdw[7];
	assign	monmdw[6] = gatead & mdw[6];
	assign	monmdw[5] = gatead & mdw[5];
	assign	monmdw[4] = gatead & mdw[4];
	assign	monmdw[3] = gatead & mdw[3];
	assign	monmdw[2] = gatead & mdw[2];
	assign	monmdw[1] = gatead & mdw[1];
	assign	monmdw[0] = gatead & mdw[0];

endmodule

/********************************************************************************/
/* K0R EVA ALU Block                                                           	*/
/*                                                          Made K.Tanaka       */
/********************************************************************************/
/* Ver1.00  New                                                                 */
/* Ver1.50  Add mem_access                            2007.05.30 K.Tanaka       */
/********************************************************************************/
module QLK0RCPUEVA0V3_ALU(
	imdr, pselcpu, pselbcd, slreg, vpa, pid, mdw, ma_pre, maw1, biten, pc, pc_inc, wdop, wdwr,
	pa_st2, pa_data_buf, pa_data_mem, pa_data_spen,
	slflash, slmirr, pc_set_brk, pc_set_dbg,
	ID_stage0, MEM_stage0, MEM_stage1,
	cpuwr, cpuwr_reg, cpurd, stage_cut, A, X, B, C, D, E, H, L, CS, ES, PSW, MAA, BCDADJ,
	A_bank0, X_bank0, B_bank0, C_bank0, D_bank0, E_bank0, H_bank0, L_bank0,
	A_bank1, X_bank1, B_bank1, C_bank1, D_bank1, E_bank1, H_bank1, L_bank1,
	A_bank2, X_bank2, B_bank2, C_bank2, D_bank2, E_bank2, H_bank2, L_bank2,
	A_bank3, X_bank3, B_bank3, C_bank3, D_bank3, E_bank3, H_bank3, L_bank3,
	A_access, X_access, B_access, C_access,
	D_access, E_access, H_access, L_access,
	INT_access, skp_block,
	intblock, PSW_block, SP_enable, CS_enable, stage_cut_br,
	buf2, buf1, buf0, SP, sp_inc, dmard, dmawr, dmawdop, waitdma,
	ivack, ivack_pre, intisp, fchiram, fchiram_skp, romrd_skp, pc_wait_flg, reg_wait,
	data_hazard_flg, data_hazard, sp_hazard,
	dec_alu_input10, dec_alu_input20,
	dec_alu_add, dec_alu_sub, dec_alu_and, dec_alu_or, dec_alu_exor,
	dec_alu_andbit, dec_alu_orbit, dec_alu_exorbit,
	dec_alu_ror, dec_alu_rol, dec_alu_shr, dec_alu_shl, dec_alu_sar,
	dec_alu_mulu, dec_alu_carry,
        dec_alu_transin, dec_alu_transout, dec_alu_bitsh, dec_alu_biten, dec_word_access,
	dec_xch_byte, dec_xchw_bc, dec_xchw_de, dec_xchw_hl,
	dec_SP_enable,
	dec_A_enable, dec_X_enable,
	dec_B_enable, dec_C_enable,
	dec_D_enable, dec_E_enable,
	dec_H_enable, dec_L_enable,
	dec_ES_enable, dec_Z_enable, dec_CY_enable, dec_AC_enable,
	dec_IE_enable, dec_ISP_enable, dec_RBS_enable,
	dec_buf0_enable, dec_buf1_enable, dec_buf2_enable,
	dec_cpuwr_enable, dec_cpurd_enable,
	dec_sp_set_enable, dec_sp_inc, dec_sp_dec,
	dec_stage_cut_brtf, dec_stage_cut_ifbr,
	dec_ifbr_not, dec_ifbr_zero, dec_ifbr_ht,
	dec_set_buf_retadr, dec_set_buf_intr,
	dec_skc, dec_sknc, dec_skz, dec_sknz, dec_skh, dec_sknh, dec_movs, dec_cmps,
	dec_ma_enable,
	skpack, skipexe, pswlock, wait_block_brtf, mem_access,
// for EVA
        SP_usr, SP_sv,
        svmod, svmodi,
        alt1, alt2,
        spinc, spdec,
        icecsgregu, icecsgrega, iceifa,
        SP0, icedo,
//
	cpuen, pswen, baseck, resb, scanmode,
	RVEON
	);

	output	[15:0]	mdw;
	output	[7:0]	biten;
	output		wdop, wdwr;
	output		cpuwr, cpuwr_reg, cpurd, stage_cut;
	output	[7:0]	A, X, B, C, D, E, H, L, buf1, buf0;
	output	[7:0]	A_bank0,X_bank0,B_bank0,C_bank0,D_bank0,E_bank0,H_bank0,L_bank0;
	output	[7:0]	A_bank1,X_bank1,B_bank1,C_bank1,D_bank1,E_bank1,H_bank1,L_bank1;
	output	[7:0]	A_bank2,X_bank2,B_bank2,C_bank2,D_bank2,E_bank2,H_bank2,L_bank2;
	output	[7:0]	A_bank3,X_bank3,B_bank3,C_bank3,D_bank3,E_bank3,H_bank3,L_bank3;
	output		A_access,X_access,B_access,C_access;
	output		D_access,E_access,H_access,L_access;
	output		INT_access;
	output	[3:0]	CS, ES, buf2;
	output		MAA;
	output	[14:0]	SP, sp_inc;
	output		skpack, skipexe;
	output	[7:0]	PSW;
	output	[1:0]	BCDADJ;
	output		skp_block;
	output		intblock;
	output		PSW_block;
	output		stage_cut_br;
	output		wait_block_brtf;
	output		mem_access;
	output		RVEON;
// for EVA
        output          spinc, spdec;
        output          SP0;
        output  [31:0]  icedo;
//

	input		SP_enable, CS_enable;
	input		pa_data_buf, pa_data_mem, pa_data_spen;
	input		pa_st2;
	input		slflash;
	input		slreg;
	input		slmirr;
	input	[15:0]	imdr;
	input		pselcpu, pselbcd;
	input	[3:0]	vpa;
	input	[31:0]	pid;
	input	[15:0]	ma_pre;
	input		maw1;
	input	[19:0]	pc, pc_inc;
	input	[7:0]	ID_stage0, MEM_stage0, MEM_stage1;
	input		dmard, dmawr, dmawdop, waitdma;
	input		ivack, ivack_pre;
	input	[1:0]	intisp;
	input		fchiram, fchiram_skp, romrd_skp;
	input		pc_wait_flg, reg_wait;
	input		pc_set_brk, pc_set_dbg;
	input		data_hazard_flg, data_hazard, sp_hazard;
	input	[3:0]	dec_alu_input10;
	input	[3:0]	dec_alu_input20;
	input	[3:0]	dec_alu_transout;
	input		dec_alu_transin;
	input	[4:0]	dec_alu_bitsh;
	input		dec_alu_biten;
	input		dec_alu_add, dec_alu_sub, dec_alu_and, dec_alu_or, dec_alu_exor;
	input		dec_alu_andbit, dec_alu_orbit, dec_alu_exorbit;
	input		dec_alu_ror, dec_alu_rol, dec_alu_shr, dec_alu_shl, dec_alu_sar;
	input		dec_alu_mulu, dec_alu_carry;
	input		dec_word_access;
	input		dec_xch_byte, dec_xchw_bc, dec_xchw_de, dec_xchw_hl;
	input		dec_SP_enable;
	input		dec_A_enable, dec_X_enable;
	input		dec_B_enable, dec_C_enable;
	input		dec_D_enable, dec_E_enable;
	input		dec_H_enable, dec_L_enable;
	input		dec_ES_enable, dec_Z_enable, dec_CY_enable, dec_AC_enable;
	input		dec_IE_enable, dec_ISP_enable, dec_RBS_enable;
	input		dec_buf0_enable, dec_buf1_enable, dec_buf2_enable;
	input		dec_cpuwr_enable, dec_cpurd_enable;
	input		dec_sp_set_enable, dec_sp_inc, dec_sp_dec;
	input		dec_stage_cut_brtf, dec_stage_cut_ifbr;
	input		dec_ifbr_not, dec_ifbr_zero, dec_ifbr_ht;
	input		dec_set_buf_retadr, dec_set_buf_intr;
	input		dec_skc, dec_sknc, dec_skz, dec_sknz, dec_skh, dec_sknh;
	input		dec_movs, dec_cmps;
	input		dec_ma_enable;
	input		pswlock;
	input		cpuen, pswen, baseck, resb;
	input		scanmode;

// for EVA
        input           svmod, svmodi;
        input           alt1, alt2;
        input           icecsgregu, icecsgrega;
        input   [2:0]   iceifa;
//

	wire	[15:0]	mdw_pre, mdw_dma;
	wire	[14:0]	sp_inc;
	wire	[15:0]	bufr;
	wire	[7:0]	PSW;
	wire	[15:0]	bitshout, exeout, muluout, aluout, aluoutpsw;
	wire		acout, cyout ,cyout1, cyout2;
	wire		PSW_enable, PSW_block_pre;
	wire		bank0, bank1, bank2, bank3;
	wire		bank_correspond;
	wire		A_access,X_access,B_access,C_access;
	wire		D_access,E_access,H_access,L_access;
	wire		wdop_pre;
	wire		sp_sfr_en;
	wire	[1:0]	bcdadj_flg;
	wire		bcdadj_low;
	wire	[1:0]	BCDADJ;
	wire	[7:0]	A_groupA,X_groupA,B_groupA,C_groupA,D_groupA,E_groupA,H_groupA,L_groupA;
	wire	[7:0]	A_groupB,X_groupB,B_groupB,C_groupB,D_groupB,E_groupB,H_groupB,L_groupB;
	wire	[7:0]	A_groupC,X_groupC,B_groupC,C_groupC,D_groupC,E_groupC,H_groupC,L_groupC;
	wire	[7:0]	MEM_stage0_groupA, MEM_stage1_groupA;
	wire	[15:0]	imdr_groupA, imdr_groupB, bufr_groupA, bufr_groupB;
	wire		cpuwr_reg;

	reg	[7:0]	biten;
// for EVA
//	reg	[14:0]	SP, sp_pre;
	reg	[14:0]	sp_pre;
//
	reg	[7:0]	A,X,B,C,D,E,H,L,buf0,buf1;
	reg	[7:0]	A_bank0,X_bank0,B_bank0,C_bank0,D_bank0,E_bank0,H_bank0,L_bank0;
	reg	[7:0]	A_bank1,X_bank1,B_bank1,C_bank1,D_bank1,E_bank1,H_bank1,L_bank1;
	reg	[7:0]	A_bank2,X_bank2,B_bank2,C_bank2,D_bank2,E_bank2,H_bank2,L_bank2;
	reg	[7:0]	A_bank3,X_bank3,B_bank3,C_bank3,D_bank3,E_bank3,H_bank3,L_bank3;
// for EVA
//	reg	[3:0]	CS,ES,buf2;
	reg	[3:0]	buf2;
//
	reg		MAA;
	reg	[1:0]	ISP;
	reg		Z,AC,CY,IE;
	reg	[1:0]	RBS;
	reg	[7:0]	aluin10, aluin11, aluin20, aluin21;
	reg	[7:0]	bitshin10, bitshin20, bitshin21;
	reg	[15:0]	transout, transin;
	reg		mem_access ;
	reg		cpuwr_pre, cpurd_pre;
	reg		fchiram_cpurd;
	reg		stage_cut, stage_cut_ifbr, stage_cut_brtf, stage_cut_alu;
	reg		wait_block_brtf;
	reg		ifbr_not, ifbr_zero, ifbr_ht;
	reg		skpack, skip_c, skip_nc, skip_z, skip_nz, skip_h, skip_nh;
	reg		intblock;
	reg		prefix_skp;
	reg	[15:0]	rdata;
	reg		PSW_block;
	reg		isp_hazard ;
	reg		sp_sfr_msk ;
	reg		RVEON;

/*------------------------------------------------------------------------------*/
/* ���̣����ϣ�									*/
/*------------------------------------------------------------------------------*/
/*   ���̣����ϣ������򤹤롣							*/
/*------------------------------------------------------------------------------*/

// �̾�MDR�Х��Υǡ�����ALU�����Ϥ��뤬��FLASH�Υǡ����꡼�ɤξ��ϡ�
// �ݻ��Хåե��˳�Ǽ���줿PID�Х��Υǡ������ɤ߽Ф���
/*------------------------------------------------------------------------------*/
/* Ver2.0  bufr(imdr)�η�ϩ��ɬ�פʻ��������Ϥ��롣				*/
/*------------------------------------------------------------------------------*/
/* Ver3.0  �ǥ��쥤�ˤ��ҥ��ɻߤ��к���ľ��(CPUV1.5���������᤹)		*/
/*------------------------------------------------------------------------------*/
	assign bufr = (pa_data_mem) ? {buf1, buf0} : imdr ;
	assign bufr_groupA = (pa_data_mem) ? {buf1, buf0} : imdr ;
	assign bufr_groupB = (pa_data_mem) ? {buf1, buf0} : imdr ;
//	assign bufr_groupA = (pa_data_mem) ? {buf1, buf0} : imdr_groupA ;
//	assign bufr_groupB = (pa_data_mem) ? {buf1, buf0} : imdr_groupB ;

// ALU���ϣ��β��̣��ӥåȤ����򤹤롣
/*------------------------------------------------------------------------------*/
/* Ver2.0  ���ѥ쥸������bufr��ɬ�פʻ���������_groupA,B,C���ѹ�		*/
/*------------------------------------------------------------------------------*/
	always @(dec_alu_input10 or vpa or A_groupB or X_groupB or B_groupB or C_groupB or D_groupB or
		E_groupB or H_groupB or L_groupB or CY or buf0 or SP or bufr_groupB) begin
		casex ({dec_alu_input10,vpa[0]})
			({4'h1,1'bx}) : aluin10 = 8'h01 ;
			({4'h3,1'bx}) : aluin10 = A_groupB ;
			({4'h4,1'bx}) : aluin10 = X_groupB ;
			({4'h5,1'bx}) : aluin10 = B_groupB ;
			({4'h6,1'bx}) : aluin10 = C_groupB ;
			({4'h7,1'bx}) : aluin10 = D_groupB ;
			({4'h8,1'bx}) : aluin10 = E_groupB ;
			({4'h9,1'bx}) : aluin10 = H_groupB ;
			({4'ha,1'bx}) : aluin10 = L_groupB ;
			({4'hb,1'bx}) : aluin10 = bufr_groupB[7:0] ;
			({4'hd,1'bx}) : aluin10 = {SP[6:0],1'b0} ;
			({4'he,1'b0}) : aluin10 = bufr_groupB[7:0] ;
			({4'he,1'b1}) : aluin10 = bufr_groupB[15:8] ;
			default : aluin10 = 8'h00 ;
		endcase
	end

// ALU���ϣ��ξ�̣��ӥåȤ����򤹤롣
/*------------------------------------------------------------------------------*/
/* Ver2.0  ���ѥ쥸������bufr��ɬ�פʻ���������_groupA,B,C���ѹ�		*/
/*------------------------------------------------------------------------------*/
	always @(dec_word_access or dec_alu_input10 or A_groupB or B_groupB or D_groupB or H_groupB or
		buf1 or SP or bufr_groupB) begin
		casex ({dec_word_access,dec_alu_input10})
			({1'b1,4'h4}) : aluin11 = A_groupB ;
			({1'b1,4'h6}) : aluin11 = B_groupB ;
			({1'b1,4'h8}) : aluin11 = D_groupB ;
			({1'b1,4'ha}) : aluin11 = H_groupB ;
			({1'b1,4'hb}) : aluin11 = bufr_groupB[15:8] ;
			({1'b1,4'hd}) : aluin11 = SP[14:7] ;
			({1'b1,4'he}) : aluin11 = bufr_groupB[15:8] ;
			default : aluin11 = 8'h00 ;
		endcase
	end

/*------------------------------------------------------------------------------*/
// Ver2.0����ή�︺�ΰ٤˥��͡��֥뿮���ɬ�פʷ�ϩ�Τߤ򳫤�
/*------------------------------------------------------------------------------*/
/* Ver3.0  ��ή�︺�θ��̤���ǧ�Ǥ��ʤ��ä�����Ver1.5���᤹			*/
/*------------------------------------------------------------------------------*/

	assign MEM_stage0_groupA = MEM_stage0 ;
	assign MEM_stage1_groupA = MEM_stage1 ;

//	assign MEM_stage0_groupA = (
//			   dec_alu_input20==4'ha	//aluin20
//			|| dec_alu_input20==4'hb	//aluin20
//			|| dec_alu_bitsh[3]		//biten,bitshin20
//			|| dec_alu_transout==4'ha	//transout[7:0]
//			|| dec_alu_shr			//bitshout
//			|| dec_alu_shl			//bitshout
//			|| dec_alu_sar			//bitshout
//			) ? MEM_stage0 : 8'h00;
//
//	assign MEM_stage1_groupA = (
//			   dec_alu_input20==4'ha	//aluin21
//			|| dec_alu_transout==4'ha	//transout[15:8]
//			) ? MEM_stage1 : 8'h00;

/*------------------------------------------------------------------------------*/
/* ���̣����ϣ�									*/
/*------------------------------------------------------------------------------*/
/*   ���̣����ϣ������򤹤롣							*/
/*------------------------------------------------------------------------------*/
/* Ver2.0  ALU��ʬ�䡣�ܡݡ��á�����						*/
/*�����������ѥ쥸������bufr��ɬ�פʻ���������_groupA,B,C���ѹ�			*/
/*------------------------------------------------------------------------------*/

// ALU���ϣ��β��̣��ӥåȤ����򤹤롣
// ADDW/SUBW SP,#byte(dec_alu_input20��5'h0b)�λ��ϥ�ɥ��������Ǥ���ʤ���
// �黻��ɬ�פʥǡ����ϥХ��ȤǤ��뤿�ᡢ��̣��ӥåȤ������̣��ӥåȤ�MEM_stage0
// �Ȥ��ä��ȹ礻����̤��Ѱդ�����
	always @(dec_alu_input20 or vpa or
		A_groupB or X_groupB or B_groupB or C_groupB or D_groupB or E_groupB or H_groupB or L_groupB or
		MEM_stage0_groupA or MEM_stage1_groupA or
		bufr_groupB or buf0 or buf2 or CY or PSW) begin
		casex ({dec_alu_input20,MEM_stage0_groupA[6:4],vpa[0]})
			({4'h1,3'hx,1'bx}) : aluin20 = 8'h01 ;
			({4'h2,3'hx,1'bx}) : aluin20 = A_groupB ;
			({4'h3,3'hx,1'bx}) : aluin20 = X_groupB ;
			({4'h4,3'hx,1'bx}) : aluin20 = B_groupB ;
			({4'h5,3'hx,1'bx}) : aluin20 = C_groupB ;
			({4'h6,3'hx,1'bx}) : aluin20 = D_groupB ;
			({4'h7,3'hx,1'bx}) : aluin20 = E_groupB ;
			({4'h8,3'hx,1'bx}) : aluin20 = H_groupB ;
			({4'h9,3'hx,1'bx}) : aluin20 = L_groupB ;
			({4'ha,3'hx,1'bx}) : aluin20 = MEM_stage0_groupA ;
			({4'hb,3'hx,1'bx}) : aluin20 = MEM_stage0_groupA ;
			({4'hc,3'hx,1'b0}) : aluin20 = bufr_groupB[7:0] ;
			({4'hc,3'hx,1'b1}) : aluin20 = bufr_groupB[15:8] ;
			({4'hd,3'hx,1'bx}) : aluin20 = {4'b0,buf2} ;
			({4'he,3'hx,1'bx}) : aluin20 = buf0 ;
			default : aluin20 = 8'h00 ;
		endcase
	end

// ALU���ϣ��ξ�̣��ӥåȤ����򤹤롣
	always @(dec_word_access or dec_alu_input20 or A_groupB or B_groupB or D_groupB or H_groupB or
		MEM_stage1_groupA or bufr_groupB or buf1 or PSW) begin
		casex ({dec_word_access,dec_alu_input20})
			({1'b1,4'h3}) : aluin21 = A_groupB ;
			({1'b1,4'h5}) : aluin21 = B_groupB ;
			({1'b1,4'h7}) : aluin21 = D_groupB ;
			({1'b1,4'h9}) : aluin21 = H_groupB ;
			({1'b1,4'ha}) : aluin21 = MEM_stage1_groupA ;
			({1'b1,4'hc}) : aluin21 = bufr_groupB[15:8] ;
			({1'b1,4'hd}) : aluin21 = PSW ;
			({1'b1,4'he}) : aluin21 = buf1 ;
			default : aluin21 = 8'h00 ;
		endcase
	end

/*------------------------------------------------------------------------------*/
/* �£ɣԣţο���								*/
/*------------------------------------------------------------------------------*/
/*   �ӥå����̿��Ǥ�ͭ���ӥåȤ���ꤹ�롣					*/
/*   dec_alu_input20 �� 0x10,0x11,0x12,0x13,0x14,0x15 �λ��ϥӥåȥ�������	*/
/*------------------------------------------------------------------------------*/
/* Ver2.0  dec_alu_bitsh �� "8,9,c,d,e,f,18,19,1c,1d" �λ��ϥӥåȥ�������      */
/*��������MEM_stage0��ɬ�פʻ���������_groupA,B,C���ѹ�				*/
/*------------------------------------------------------------------------------*/

// �ӥå����̿��Ǥʤ��������ӥåȤˣ���Ω�Ƥ롣
	always @(dec_alu_biten or MEM_stage0) begin
		if (dec_alu_biten == 1'b1) begin
			casex (MEM_stage0[6:4])
				3'h1 : biten = 8'b0000_0010 ;
				3'h2 : biten = 8'b0000_0100 ;
				3'h3 : biten = 8'b0000_1000 ;
				3'h4 : biten = 8'b0001_0000 ;
				3'h5 : biten = 8'b0010_0000 ;
				3'h6 : biten = 8'b0100_0000 ;
				3'h7 : biten = 8'b1000_0000 ;
				default : biten = 8'b0000_0001 ;
			endcase
		end
		else biten = 8'b1111_1111 ;
	end

/*------------------------------------------------------------------------------*/
/* ���̣ձ黻									*/
/*------------------------------------------------------------------------------*/
/*   ���̣ձ黻�μ�������򤹤롣						*/
/*------------------------------------------------------------------------------*/
/* Ver2.0  MEM_stage0��ɬ�פʻ���������_groupA,B,C���ѹ�			*/
/*------------------------------------------------------------------------------*/

// �黻��¹Ԥ��륿���ߥ󥰥ѥ��Ȥ���ʳ��Υѥ�����̤���٤˳��ز����롣
	QLK0RCPUEVA0V3_EXE exe (.aluin10(aluin10), .aluin11(aluin11), .aluin20(aluin20), .aluin21(aluin21), .CY(CY),
			     .dec_alu_add(dec_alu_add), .dec_alu_sub(dec_alu_sub), .dec_alu_and(dec_alu_and), 
			     .dec_alu_or(dec_alu_or), .dec_alu_exor(dec_alu_exor), 
			     .dec_alu_carry(dec_alu_carry), .dec_word_access(dec_word_access),
			     .exeout(exeout), .acout(acout), .cyout(cyout1) );

/*------------------------------------------------------------------------------*/
/* Ver2.0  ALU��ʬ�䡣�軻������						*/
/*------------------------------------------------------------------------------*/

	assign muluout = (dec_alu_mulu) ? (A_groupB * X_groupB) : 16'h0000;

/*------------------------------------------------------------------------------*/
/* Ver2.0  ALU��ʬ�䡣ž���Υ��ꥢ��������������				*/
/*------------------------------------------------------------------------------*/

	always @(dec_alu_transout or vpa or A_groupA or X_groupA or B_groupA or C_groupA or D_groupA or
		E_groupA or H_groupA or L_groupA or MEM_stage0_groupA or buf0 or buf2) begin
		casex ({dec_alu_transout,vpa[0]})
			({4'h1,1'bx}) : transout[7:0] = 8'h01 ;
			({4'h2,1'bx}) : transout[7:0] = A_groupA ;
			({4'h3,1'bx}) : transout[7:0] = X_groupA ;
			({4'h4,1'bx}) : transout[7:0] = B_groupA ;
			({4'h5,1'bx}) : transout[7:0] = C_groupA ;
			({4'h6,1'bx}) : transout[7:0] = D_groupA ;
			({4'h7,1'bx}) : transout[7:0] = E_groupA ;
			({4'h8,1'bx}) : transout[7:0] = H_groupA ;
			({4'h9,1'bx}) : transout[7:0] = L_groupA ;
			({4'ha,1'bx}) : transout[7:0] = MEM_stage0_groupA ;
			({4'hd,1'bx}) : transout[7:0] = {4'b0,buf2} ;
			({4'he,1'bx}) : transout[7:0] = buf0 ;
			default : transout[7:0] = 8'h00 ;
		endcase
	end
	always @(dec_word_access or dec_alu_transout or A_groupA or B_groupA or D_groupA or H_groupA or
		MEM_stage1_groupA or PSW or buf1) begin
		casex ({dec_word_access,dec_alu_transout})
			({1'b1,4'h3}) : transout[15:8] = A_groupA ;
			({1'b1,4'h5}) : transout[15:8] = B_groupA ;
			({1'b1,4'h7}) : transout[15:8] = D_groupA ;
			({1'b1,4'h9}) : transout[15:8] = H_groupA ;
			({1'b1,4'ha}) : transout[15:8] = MEM_stage1_groupA ;
			({1'b1,4'hd}) : transout[15:8] = PSW ;
			({1'b1,4'he}) : transout[15:8] = buf1 ;
			({1'b1,4'hf}) : transout[15:8] = PSW ;
			default : transout[15:8] = 8'h00 ;
		endcase
	end

/*------------------------------------------------------------------------------*/
/* Ver2.0  ALU��ʬ�䡣ž���Υ��꤫�����������				*/
/*------------------------------------------------------------------------------*/

	always @(dec_alu_transin or vpa or bufr_groupA) begin
		casex ({dec_alu_transin,vpa[0]})
			({1'b1,1'b0}) : transin[7:0] = bufr_groupA[7:0] ;
			({1'b1,1'b1}) : transin[7:0] = bufr_groupA[15:8] ;
			default : transin[7:0] = 8'h00 ;
		endcase
	end
	always @(dec_word_access or dec_alu_transin or bufr_groupA) begin
		casex ({dec_word_access,dec_alu_transin})
			({1'b1,1'b1}) : transin[15:8] = bufr_groupA[15:8] ;
			default : transin[15:8] = 8'h00 ;
		endcase
	end

/*------------------------------------------------------------------------------*/
/* Ver2.0  ALU��ʬ�䡣���եȡ��ӥå�̿������					*/
/*------------------------------------------------------------------------------*/

// ALU����1�β��̣��ӥåȤ����򤹤롣

        always @(dec_alu_bitsh or vpa or A_groupB or bufr_groupB or CY) begin
                casex ({dec_alu_bitsh, vpa[0]})
                        ({5'b1100x,1'bx}) : bitshin10 = 8'h01 ;
                        ({5'b1110x,1'bx}) : bitshin10 = A_groupB ;
                        ({5'b0110x,1'b0}) : bitshin10 = bufr_groupB[7:0] ;
                        ({5'b0110x,1'b1}) : bitshin10 = bufr_groupB[15:8] ;
                        ({5'b0100x,1'bx}) : bitshin10 = {7'h00,CY} ;
                        ({5'b10001,1'bx}) : bitshin10 = {7'h00,CY} ;
                        default : bitshin10 = 8'h00 ;
                endcase
        end

// ALU���ϣ��β��̣��ӥåȤ����򤹤롣
        always @(dec_alu_bitsh or vpa or A_groupB or X_groupB or B_groupB or C_groupB or
                MEM_stage0_groupA or bufr_groupB or CY) begin
                casex ({dec_alu_bitsh, MEM_stage0_groupA[6:4], vpa[0]})
                        ({5'bx0001,3'hx,1'bx}) : bitshin20 = 8'hff ;			// 0x01, 0x11
                        ({5'b00010,3'hx,1'bx}) : bitshin20 = A_groupB ;			// 0x02
                        ({5'b00011,3'hx,1'bx}) : bitshin20 = X_groupB ;			// 0x03
                        ({5'b00100,3'hx,1'bx}) : bitshin20 = B_groupB ;			// 0x04
                        ({5'b00101,3'hx,1'bx}) : bitshin20 = C_groupB ;			// 0x05
                        ({5'bx1000,3'h0,1'b0}) : bitshin20 = {7'b0,bufr_groupB[0]} ;	// 0x08, 0x18
                        ({5'bx1000,3'h1,1'b0}) : bitshin20 = {7'b0,bufr_groupB[1]} ;	// 0x08, 0x18
                        ({5'bx1000,3'h2,1'b0}) : bitshin20 = {7'b0,bufr_groupB[2]} ;	// 0x08, 0x18
                        ({5'bx1000,3'h3,1'b0}) : bitshin20 = {7'b0,bufr_groupB[3]} ;	// 0x08, 0x18
                        ({5'bx1000,3'h4,1'b0}) : bitshin20 = {7'b0,bufr_groupB[4]} ;	// 0x08, 0x18
                        ({5'bx1000,3'h5,1'b0}) : bitshin20 = {7'b0,bufr_groupB[5]} ;	// 0x08, 0x18
                        ({5'bx1000,3'h6,1'b0}) : bitshin20 = {7'b0,bufr_groupB[6]} ;	// 0x08, 0x18
                        ({5'bx1000,3'h7,1'b0}) : bitshin20 = {7'b0,bufr_groupB[7]} ;	// 0x08, 0x18
                        ({5'bx1000,3'h0,1'b1}) : bitshin20 = {7'b0,bufr_groupB[8]} ;	// 0x08, 0x18
                        ({5'bx1000,3'h1,1'b1}) : bitshin20 = {7'b0,bufr_groupB[9]} ;	// 0x08, 0x18
                        ({5'bx1000,3'h2,1'b1}) : bitshin20 = {7'b0,bufr_groupB[10]} ;	// 0x08, 0x18
                        ({5'bx1000,3'h3,1'b1}) : bitshin20 = {7'b0,bufr_groupB[11]} ;	// 0x08, 0x18
                        ({5'bx1000,3'h4,1'b1}) : bitshin20 = {7'b0,bufr_groupB[12]} ;	// 0x08, 0x18
                        ({5'bx1000,3'h5,1'b1}) : bitshin20 = {7'b0,bufr_groupB[13]} ;	// 0x08, 0x18
                        ({5'bx1000,3'h6,1'b1}) : bitshin20 = {7'b0,bufr_groupB[14]} ;	// 0x08, 0x18
                        ({5'bx1000,3'h7,1'b1}) : bitshin20 = {7'b0,bufr_groupB[15]} ;	// 0x08, 0x18
                        ({5'bx1001,3'h0,1'bx}) : bitshin20 = {7'b0,A_groupB[0]} ;	// 0x09, 0x19
                        ({5'bx1001,3'h1,1'bx}) : bitshin20 = {7'b0,A_groupB[1]} ;	// 0x09, 0x19
                        ({5'bx1001,3'h2,1'bx}) : bitshin20 = {7'b0,A_groupB[2]} ;	// 0x09, 0x19
                        ({5'bx1001,3'h3,1'bx}) : bitshin20 = {7'b0,A_groupB[3]} ;	// 0x09, 0x19
                        ({5'bx1001,3'h4,1'bx}) : bitshin20 = {7'b0,A_groupB[4]} ;	// 0x09, 0x19
                        ({5'bx1001,3'h5,1'bx}) : bitshin20 = {7'b0,A_groupB[5]} ;	// 0x09, 0x19
                        ({5'bx1001,3'h6,1'bx}) : bitshin20 = {7'b0,A_groupB[6]} ;	// 0x09, 0x19
                        ({5'bx1001,3'h7,1'bx}) : bitshin20 = {7'b0,A_groupB[7]} ;	// 0x09, 0x19
                        ({5'b01110,3'h0,1'b0}) : bitshin20 = {bufr_groupB[7:1],CY} ;	// 0x0e
                        ({5'b01110,3'h1,1'b0}) : bitshin20 = {bufr_groupB[7:2],CY,bufr_groupB[0]} ;	// 0x0e
                        ({5'b01110,3'h2,1'b0}) : bitshin20 = {bufr_groupB[7:3],CY,bufr_groupB[1:0]} ;	// 0x0e
                        ({5'b01110,3'h3,1'b0}) : bitshin20 = {bufr_groupB[7:4],CY,bufr_groupB[2:0]} ;	// 0x0e
                        ({5'b01110,3'h4,1'b0}) : bitshin20 = {bufr_groupB[7:5],CY,bufr_groupB[3:0]} ;	// 0x0e
                        ({5'b01110,3'h5,1'b0}) : bitshin20 = {bufr_groupB[7:6],CY,bufr_groupB[4:0]} ;	// 0x0e
                        ({5'b01110,3'h6,1'b0}) : bitshin20 = {bufr_groupB[7],CY,bufr_groupB[5:0]} ;	// 0x0e
                        ({5'b01110,3'h7,1'b0}) : bitshin20 = {CY,bufr_groupB[6:0]} ;	// 0x0e
                        ({5'b01110,3'h0,1'b1}) : bitshin20 = {bufr_groupB[15:9],CY} ;	// 0x0e
                        ({5'b01110,3'h1,1'b1}) : bitshin20 = {bufr_groupB[15:10],CY,bufr_groupB[8]} ;	// 0x0e
                        ({5'b01110,3'h2,1'b1}) : bitshin20 = {bufr_groupB[15:11],CY,bufr_groupB[9:8]} ;	// 0x0e
                        ({5'b01110,3'h3,1'b1}) : bitshin20 = {bufr_groupB[15:12],CY,bufr_groupB[10:8]} ;// 0x0e
                        ({5'b01110,3'h4,1'b1}) : bitshin20 = {bufr_groupB[15:13],CY,bufr_groupB[11:8]} ;// 0x0e
                        ({5'b01110,3'h5,1'b1}) : bitshin20 = {bufr_groupB[15:14],CY,bufr_groupB[12:8]} ;// 0x0e
                        ({5'b01110,3'h6,1'b1}) : bitshin20 = {bufr_groupB[15],CY,bufr_groupB[13:8]} ;	// 0x0e
                        ({5'b01110,3'h7,1'b1}) : bitshin20 = {CY,bufr_groupB[14:8]} ;	// 0x0e
                        ({5'bx1101,3'h0,1'bx}) : bitshin20 = 8'h01 ;			// 0x0d, 0x1d
                        ({5'bx1101,3'h1,1'bx}) : bitshin20 = 8'h02 ;			// 0x0d, 0x1d
                        ({5'bx1101,3'h2,1'bx}) : bitshin20 = 8'h04 ;			// 0x0d, 0x1d
                        ({5'bx1101,3'h3,1'bx}) : bitshin20 = 8'h08 ;			// 0x0d, 0x1d
                        ({5'bx1101,3'h4,1'bx}) : bitshin20 = 8'h10 ;			// 0x0d, 0x1d
                        ({5'bx1101,3'h5,1'bx}) : bitshin20 = 8'h20 ;			// 0x0d, 0x1d
                        ({5'bx1101,3'h6,1'bx}) : bitshin20 = 8'h40 ;			// 0x0d, 0x1d
                        ({5'bx1101,3'h7,1'bx}) : bitshin20 = 8'h80 ;			// 0x0d, 0x1d
                        ({5'bx1100,3'h0,1'bx}) : bitshin20 = 8'hfe ;			// 0x0c, 0x1c
                        ({5'bx1100,3'h1,1'bx}) : bitshin20 = 8'hfd ;			// 0x0c, 0x1c
                        ({5'bx1100,3'h2,1'bx}) : bitshin20 = 8'hfb ;			// 0x0c, 0x1c
                        ({5'bx1100,3'h3,1'bx}) : bitshin20 = 8'hf7 ;			// 0x0c, 0x1c
                        ({5'bx1100,3'h4,1'bx}) : bitshin20 = 8'hef ;			// 0x0c, 0x1c
                        ({5'bx1100,3'h5,1'bx}) : bitshin20 = 8'hdf ;			// 0x0c, 0x1c
                        ({5'bx1100,3'h6,1'bx}) : bitshin20 = 8'hbf ;			// 0x0c, 0x1c
                        ({5'bx1100,3'h7,1'bx}) : bitshin20 = 8'h7f ;			// 0x0c, 0x1c
                        ({5'b01111,3'h0,1'bx}) : bitshin20 = {A_groupB[7:1],CY} ;		// 0x0f
                        ({5'b01111,3'h1,1'bx}) : bitshin20 = {A_groupB[7:2],CY,A_groupB[0]} ;	// 0x0f
                        ({5'b01111,3'h2,1'bx}) : bitshin20 = {A_groupB[7:3],CY,A_groupB[1:0]} ;	// 0x0f
                        ({5'b01111,3'h3,1'bx}) : bitshin20 = {A_groupB[7:4],CY,A_groupB[2:0]} ;	// 0x0f
                        ({5'b01111,3'h4,1'bx}) : bitshin20 = {A_groupB[7:5],CY,A_groupB[3:0]} ;	// 0x0f
                        ({5'b01111,3'h5,1'bx}) : bitshin20 = {A_groupB[7:6],CY,A_groupB[4:0]} ;	// 0x0f
                        ({5'b01111,3'h6,1'bx}) : bitshin20 = {A_groupB[7],CY,A_groupB[5:0]} ;	// 0x0f
                        ({5'b01111,3'h7,1'bx}) : bitshin20 = {CY,A_groupB[6:0]} ;		// 0x0f
                        default : bitshin20 = 8'h00 ;
                endcase
        end

// ALU���ϣ��ξ�̣��ӥåȤ����򤹤롣
        always @(dec_word_access or dec_alu_bitsh or A_groupB or B_groupB ) begin
                casex ({dec_word_access,dec_alu_bitsh })
                        ({1'b1,5'h03}) : bitshin21 = A_groupB ;
                        ({1'b1,5'h05}) : bitshin21 = B_groupB ;
                        default : bitshin21 = 8'h00 ;
                endcase
        end

/*------------------------------------------------------------------------------*/
/* ���̣ձ黻2                                                                  */
/*------------------------------------------------------------------------------*/

// �黻��¹Ԥ��륿���ߥ󥰥ѥ��Ȥ���ʳ��Υѥ�����̤���٤˳��ز����롣
        QLK0RCPUEVA0V3_EXE2 exe2 (.bitshin10(bitshin10), .bitshin20(bitshin20), .bitshin21(bitshin21), .CY(CY),
                               .dec_alu_andbit(dec_alu_andbit), .dec_alu_orbit(dec_alu_orbit), 
		  	       .dec_alu_exorbit(dec_alu_exorbit), .dec_alu_ror(dec_alu_ror),
                               .dec_alu_rol(dec_alu_rol), .dec_alu_shr(dec_alu_shr), .dec_alu_shl(dec_alu_shl),
                               .dec_alu_sar(dec_alu_sar), .dec_alu_carry(dec_alu_carry),
                               .MEM_stage0h(MEM_stage0_groupA[7:4]), .dec_word_access(dec_word_access),
                               .bitshout(bitshout), .cyout(cyout2) );

/*------------------------------------------------------------------------------*/
/* Ver2.0��ALU�α黻���							*/
/*------------------------------------------------------------------------------*/
/*   aluoutpsw:PSW�α黻�˻��Ѥ��롣			 			*/
/*   aluout   :�黻��̤˻��Ѥ��롣			 			*/
/*------------------------------------------------------------------------------*/

	assign aluout = exeout | transout | transin | muluout | bitshout ;
	assign aluoutpsw = exeout | bitshout ;
	assign cyout  = cyout1 | cyout2 ;

/*------------------------------------------------------------------------------*/
/* ����ե饰�쥸���� ��							*/
/*------------------------------------------------------------------------------*/
/*   ���̣ս��Ϥ����λ����åȤ���롣						*/
/*   �Уӣפ˴ޤޤ�롣								*/
/*------------------------------------------------------------------------------*/
/* Ver2.0��aluout��aluoutpsw���ѹ�						*/
/*��������aluoutpsw���ѹ������ݤ�dec_movs�λ���aluoutpsw�˥ǡ������ΤäƤ��ʤ�	*/
/*���������١�ľ��X�쥸�������ͤ�Ƚ�ꤹ�롣					*/
/*------------------------------------------------------------------------------*/

// ������������ȯ�������ݻ�����롣
// �ǥ���������PSW�����򤵤줿���ALU���Ϥ����ꡢľ�ܥ��ꥢ�����������ä����MDW�����롣
// INT�������ˤ�볰���������ȤǤ�PSW�ϥ������Ȥ��ʤ���
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) Z <= 1'b0 ;
		else if (cpuen || pswen) begin
			if (reg_wait || pswlock) Z <= Z ;
			else if (PSW_enable) Z <= aluoutpsw[14] ;
			else if (dec_Z_enable) begin
				if      (dec_word_access && aluoutpsw == 16'h0000) Z <= 1'b1 ;
				else if (!dec_word_access && aluoutpsw[7:0] == 8'h00) Z <= 1'b1 ;
				else Z <= 1'b0 ;
			end
			else if (dec_movs) begin
				if (X_groupB == 8'h00) Z <= 1'b1 ;
				else Z <= 1'b0 ;
			end
			else if (pselcpu && cpuwr) begin
				casex (vpa)
					4'ha : Z <= mdw_pre[6] ;
					default	: Z <= Z ;
				endcase
			end
		end
	end

/*------------------------------------------------------------------------------*/
/* ����꡼�ե饰�쥸���� �ã�							*/
/*------------------------------------------------------------------------------*/
/*   ���̣դα黻�ǥ���꡼��ȯ��������祻�åȤ���롣				*/
/*   �Уӣפ˴ޤޤ�롣								*/
/*   dec_alu_input20 �� 0x10,0x11,0x12,0x13,0x14,0x15 �λ��ϥӥåȥ�������	*/
/*------------------------------------------------------------------------------*/
/* Ver2.0 aluout��aluoutpsw���ѹ�						*/
/*�����������ѥ쥸������ɬ�פʻ���������_groupA,B,C���ѹ�			*/
/*��������dec_alu_bitsh = 0x08,0x09,0x01,0x11 && dec_CY_enable = 1		*/
/*��������						-> CY = aluoutpsw[0]	*/
/*------------------------------------------------------------------------------*/

// ������������ȯ�������ݻ�����롣
// �ǥ���������PSW�����򤵤줿���ALU���Ϥ����ꡢľ�ܥ��ꥢ�����������ä����MDW�����롣
// INT�������ˤ�볰���������ȤǤ�PSW�ϥ������Ȥ��ʤ���
// ADDC/SUBC̿��ǡ��ϥ����ɤ�ȯ��������硢�����ʱ黻��̤�CY������ʤ��Ѥˡ�data_hazard������ݻ����롣
// cyout����������BCDADJ�쥸���������򤵤�Ƥ���С�CY�Ȥ�OR���롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) CY <= 1'b0 ;
		else if (cpuen || pswen) begin
			if (reg_wait || data_hazard || pswlock) CY <= CY ;
			else if (PSW_enable) CY <= aluoutpsw[8] ;
			else if (dec_movs) CY <= (A_groupB == 8'h00) | (X_groupB == 8'h00) ;
			else if (dec_CY_enable) begin
				if ((dec_alu_bitsh == 5'h01)|(dec_alu_bitsh == 5'h08)|(dec_alu_bitsh == 5'h09)|(dec_alu_bitsh == 5'h11)) CY <= aluoutpsw[0] ;
				else if (dec_cmps) CY <= (aluoutpsw[7:0] != 8'h00) | (A_groupB == 8'h00) | (aluin10 == 8'h00) ;
				else CY <= cyout | (CY & pselbcd) ;
			end
			else if (pselcpu && cpuwr) begin
				casex (vpa)
					4'ha : CY <= mdw_pre[0] ;
					default	: CY <= CY ;
				endcase
			end
		end
	end

/*------------------------------------------------------------------------------*/
/* �������꡼�ե饰�쥸���� ����						*/
/*------------------------------------------------------------------------------*/
/*   ���̣ձ黻���������꡼��ȯ��������祻�åȤ���롣			*/
/*   �Уӣפ˴ޤޤ�롣								*/
/*------------------------------------------------------------------------------*/
/* Ver2.0 aluout��aluoutpsw���ѹ�						*/
/*------------------------------------------------------------------------------*/

// ������������ȯ�������ݻ�����롣
// �ǥ���������PSW�����򤵤줿���ALU���Ϥ����ꡢľ�ܥ��ꥢ�����������ä����MDW�����롣
// INT�������ˤ�볰���������ȤǤ�PSW�ϥ������Ȥ��ʤ���
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) AC <= 1'b0 ;
		else if (cpuen || pswen) begin
			if (reg_wait || pswlock) AC <= AC ;
			else if (PSW_enable) AC <= aluoutpsw[12] ;
			else if (dec_AC_enable) AC <= acout ;
			else if (pselcpu && cpuwr) begin
				casex (vpa)
					4'ha : AC <= mdw_pre[4] ;
					default	: AC <= AC ;
				endcase
			end
		end
	end

/*------------------------------------------------------------------------------*/
/* �����ߵ��ĥե饰�쥸���� �ɣ�						*/
/*------------------------------------------------------------------------------*/
/*   �����߼����դ���Ƚ�ꤹ�롣						*/
/*   �Уӣפ˴ޤޤ�롣								*/
/*------------------------------------------------------------------------------*/
/* Ver2.0 aluout��aluoutpsw���ѹ�						*/
/*------------------------------------------------------------------------------*/

// ������������ȯ�������ݻ�����롣
// �ǥ���������PSW�����򤵤줿���ALU���Ϥ����ꡢľ�ܥ��ꥢ�����������ä����MDW�����롣
// INT�������ˤ�볰���������ȤǤ�PSW�ϥ������Ȥ��ʤ���
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) IE <= 1'b0 ;
		else if (cpuen || pswen) begin
			if (reg_wait || pswlock) IE <= IE ;
			else if (PSW_enable) IE <= aluoutpsw[15] ;
			else if (dec_IE_enable) IE <= aluoutpsw[0] ;
			else if (pc_set_brk | pc_set_dbg) IE <= 1'b0 ;
			else if (pselcpu && cpuwr) begin
				casex (vpa)
					4'ha : IE <= mdw_pre[7] ;
					default	: IE <= IE ;
				endcase
			end
		end
	end

/*------------------------------------------------------------------------------*/
/* �쥸�����Х�����ե饰�쥸���� �ң£�					*/
/*------------------------------------------------------------------------------*/
/*   �쥸�����Х󥯤򼨤���							*/
/*   �Уӣפ˴ޤޤ�롣                                                         */
/*------------------------------------------------------------------------------*/
/* Ver2.0 aluout��aluoutpsw���ѹ�						*/
/*------------------------------------------------------------------------------*/

// ������������ȯ�������ݻ�����롣
// �ǥ���������PSW�����򤵤줿���ALU���Ϥ����ꡢľ�ܥ��ꥢ�����������ä����MDW�����롣
// SEL̿��ϥ��ڥ�������˥Х󥯤������ޤ�Ƥ���Τǡ�
// �¹Ի���ALU���̤���MEM���ơ����Υǡ��������롣
// INT�������ˤ�볰���������ȤǤ�PSW�ϥ������Ȥ��ʤ���
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) RBS <= 2'b0 ;
		else if (cpuen || pswen) begin
			if (reg_wait || pswlock) RBS <= RBS ;
			else if (PSW_enable) RBS <= {aluoutpsw[13],aluoutpsw[11]} ;
			else if (dec_RBS_enable) begin
				if (dec_alu_input20 == 4'ha) RBS <= aluoutpsw[5:4] ;
				else RBS <= {aluoutpsw[5],aluoutpsw[3]} ;
			end
			else if (pselcpu && cpuwr) begin
				casex (vpa)
					4'ha : RBS <= {mdw_pre[5],mdw_pre[3]} ;
					default	: RBS <= RBS ;
				endcase
			end
		end
	end

/*------------------------------------------------------------------------------*/
/* ������ͥ���̥ե饰�쥸���� �ɣӣ�					*/
/*------------------------------------------------------------------------------*/
/*   �����ߤ�ͥ���̤򼨤���							*/
/*   �Уӣפ˴ޤޤ�롣								*/
/*------------------------------------------------------------------------------*/

// �����߼¹Ի��˥ϥ����ɤ�ȯ���������ˣ��Ȥʤ롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) isp_hazard <= 1'b0 ;
		else if (cpuen) begin
			if (data_hazard && ivack) isp_hazard <= 1'b1 ;
			else isp_hazard <= 1'b0 ;
		end
	end

// ������������ȯ�����ȳ����߼¹Ի��Υϥ����ɤ��ݻ�����롣
// ������ȯ�������̾�ivack_pre��ISP�򹹿����뤬��
// �����߼¹Ի��˥ϥ����ɤ�ȯ����������isp_hazard�ǹ������롣
// INT�������ˤ�볰���������ȤǤ�PSW�ϥ������Ȥ��ʤ���
/*------------------------------------------------------------------------------*/
/* Ver2.0 aluout��aluoutpsw���ѹ�						*/
/*------------------------------------------------------------------------------*/

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) ISP <= 2'b11 ;
		else if (cpuen || pswen) begin
			if (reg_wait || (data_hazard && ivack) || pswlock) ISP <= ISP ;
			else if (PSW_enable) ISP <= {aluoutpsw[10],aluoutpsw[9]} ;
			else if (ivack_pre || isp_hazard) ISP <= intisp ;
			else if (dec_ISP_enable) ISP <= aluoutpsw[2:1] ;
			else if (pselcpu && cpuwr) begin
				casex (vpa)
					4'ha : ISP <= mdw_pre[2:1] ;
					default	: ISP <= ISP ;
				endcase
			end
		end
	end

/*------------------------------------------------------------------------------*/
/* �ץ���ॹ�ơ�������� �Уӣ�						*/
/*------------------------------------------------------------------------------*/
/*   �ɣš��ڡ��ң£ӣ������á��ң£ӣ����ɣӣС��ã٤ǹ�������롣		*/
/*------------------------------------------------------------------------------*/

// �ץ���ॹ�ơ��������
	assign PSW = {IE,Z,RBS[1],AC,RBS[0],ISP,CY} ;

// PSW���򿮹档�ǥ���������PSW�����򤵤줿��磱�Ȥʤ롣
	assign PSW_enable = dec_IE_enable & dec_Z_enable & dec_RBS_enable & dec_AC_enable & dec_ISP_enable & dec_CY_enable ;

// PSW�˥��������������ˣ��Ȥʤ롣INT�ޥ����IF/MK�쥸�����ؤΥ��������ȹ�碌�ơ�
// �����������ȿ���Ȥʤ롣
	assign INT_access = dec_IE_enable | PSW_enable ;

// PSW�ؤΥ��ꥢ��������ȼ�����ʬ��̿�᤬�¹Ԥ��줿��磱�Ȥʤ롣
	assign PSW_block_pre = pselcpu & (vpa == 4'ha) & dec_stage_cut_brtf ;

// ��������α�װ���PSW�ؤΥ��ꥢ��������ȼ�����ʬ��̿�᤬�¹Ԥ��줿��磱�Ȥʤ롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) PSW_block <= 1'b0 ;
		else if (cpuen) begin
			if (reg_wait)	PSW_block <= PSW_block ;
			else		PSW_block <= PSW_block_pre ;
		end
	end

// ��������α�װ���PSW��������磱�Ȥʤ롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) intblock <= 1'b0 ;
		else if (cpuen) begin
			if (reg_wait)	intblock <= intblock ;
			else		intblock <= PSW_enable ;
		end
	end

/*------------------------------------------------------------------------------*/
/* Ver3.0									*/
/* ����������߼�������쥸���� RVEON						*/
/*------------------------------------------------------------------------------*/
	always @(posedge baseck or negedge resb) begin
		if (!resb) 	RVEON <= 1'b0 ;
		else if (cpuen) begin
			if (reg_wait)	RVEON <= RVEON ;
			else if (pselbcd & cpuwr) begin
				casex ({vpa}) 
					(4'hF) : RVEON <= mdw_pre[8] ;
					default : RVEON <= RVEON ;
				endcase
			end
		end
	end
/*------------------------------------------------------------------------------*/
/* ���ѥ쥸����									*/
/*------------------------------------------------------------------------------*/
/*   ���Х��ȤΣ����ء��¡��á��ġ��š��ȡ��̥쥸�����ߣ��Х󥯤ǹ�������롣	*/
/*------------------------------------------------------------------------------*/

// for EVA

        reg     [31:0]  icedo;
        reg     [7:0]   A_sv, X_sv, B_sv, C_sv, D_sv, E_sv, H_sv, L_sv;

        always @(icecsgregu or icecsgrega or iceifa or
                 A_sv or X_sv or B_sv or C_sv or D_sv or E_sv or H_sv or L_sv or
                 A_bank0 or X_bank0 or B_bank0 or C_bank0 or D_bank0 or E_bank0 or H_bank0 or L_bank0 or
                 A_bank1 or X_bank1 or B_bank1 or C_bank1 or D_bank1 or E_bank1 or H_bank1 or L_bank1 or
                 A_bank2 or X_bank2 or B_bank2 or C_bank2 or D_bank2 or E_bank2 or H_bank2 or L_bank2 or
                 A_bank3 or X_bank3 or B_bank3 or C_bank3 or D_bank3 or E_bank3 or H_bank3 or L_bank3 ) begin
                casex ({icecsgregu,icecsgrega,iceifa})
                        5'b10_111 : icedo = {H_bank0,L_bank0,D_bank0,E_bank0} ;
                        5'b10_110 : icedo = {B_bank0,C_bank0,A_bank0,X_bank0} ;
                        5'b10_101 : icedo = {H_bank1,L_bank1,D_bank1,E_bank1} ;
                        5'b10_100 : icedo = {B_bank1,C_bank1,A_bank1,X_bank1} ;
                        5'b10_011 : icedo = {H_bank2,L_bank2,D_bank2,E_bank2} ;
                        5'b10_010 : icedo = {B_bank2,C_bank2,A_bank2,X_bank2} ;
                        5'b10_001 : icedo = {H_bank3,L_bank3,D_bank3,E_bank3} ;
                        5'b10_000 : icedo = {B_bank3,C_bank3,A_bank3,X_bank3} ;
                        5'b01_xx1 : icedo = {H_sv,L_sv,D_sv,E_sv} ;
                        5'b01_xx0 : icedo = {B_sv,C_sv,A_sv,X_sv} ;
                        5'b00_xxx : icedo = 32'b0 ;
                        default : icedo = 32'b0 ;
                endcase
        end

        wire sel_svmod_reg = svmod & ~alt2 ;
//

// RBS���ͤ˱����Ƴ�������Х󥯿��椬���Ȥʤ롣
	assign bank0 = (RBS == 2'h0) ;
	assign bank1 = (RBS == 2'h1) ;
	assign bank2 = (RBS == 2'h2) ;
	assign bank3 = (RBS == 2'h3) ;

// RBS���ͤ˱����Ƴƥ쥸�����ΥХ󥯤����򤹤롣
	always @(RBS or
// for EVA
                 sel_svmod_reg or A_sv or X_sv or B_sv or C_sv or D_sv or E_sv or H_sv or L_sv or
//
		 A_bank0 or X_bank0 or B_bank0 or C_bank0 or D_bank0 or E_bank0 or H_bank0 or L_bank0 or
		 A_bank1 or X_bank1 or B_bank1 or C_bank1 or D_bank1 or E_bank1 or H_bank1 or L_bank1 or
		 A_bank2 or X_bank2 or B_bank2 or C_bank2 or D_bank2 or E_bank2 or H_bank2 or L_bank2 or
		 A_bank3 or X_bank3 or B_bank3 or C_bank3 or D_bank3 or E_bank3 or H_bank3 or L_bank3 ) begin
// for EVA
                if (sel_svmod_reg) begin
                                {A,X,B,C,D,E,H,L} = {A_sv,X_sv,B_sv,C_sv,D_sv,E_sv,H_sv,L_sv} ;
                end
                else begin
//
		case (RBS)
			2'b00 : {A,X,B,C,D,E,H,L} = {A_bank0,X_bank0,B_bank0,C_bank0,D_bank0,E_bank0,H_bank0,L_bank0} ;
			2'b01 : {A,X,B,C,D,E,H,L} = {A_bank1,X_bank1,B_bank1,C_bank1,D_bank1,E_bank1,H_bank1,L_bank1} ;
			2'b10 : {A,X,B,C,D,E,H,L} = {A_bank2,X_bank2,B_bank2,C_bank2,D_bank2,E_bank2,H_bank2,L_bank2} ;
			2'b11 : {A,X,B,C,D,E,H,L} = {A_bank3,X_bank3,B_bank3,C_bank3,D_bank3,E_bank3,H_bank3,L_bank3} ;
		endcase
// for EVA
		end
//
	end

/*------------------------------------------------------------------------------*/
/* Ver2.0 ��ή�︺�ΰ٤˥��͡��֥뿮���ɬ�פʷ�ϩ�Τߤ򳫤�			*/
/*------------------------------------------------------------------------------*/
/* Ver3.0 ��ή�︺�θ��̤���ǧ�Ǥ��ʤ��ä�����Ver1.5���᤹			*/
/*------------------------------------------------------------------------------*/

	assign A_groupA = A;
	assign A_groupB = A;
	assign A_groupC = A;
	assign X_groupA = X;
	assign X_groupB = X;
	assign X_groupC = X;
	assign B_groupA = B;
	assign B_groupB = B;
	assign B_groupC = B;
	assign C_groupA = C;
	assign C_groupB = C;
	assign C_groupC = C;
	assign D_groupA = D;
	assign D_groupB = D;
	assign D_groupC = D;
	assign E_groupA = E;
	assign E_groupB = E;
	assign E_groupC = E;
	assign H_groupA = H;
	assign H_groupB = H;
	assign H_groupC = H;
	assign L_groupA = L;
	assign L_groupB = L;
	assign L_groupC = L;
//	assign imdr_groupA = imdr;
	assign imdr_groupB = imdr;

//	assign A_groupA = (dec_alu_transout==4'h2		//transout[7:0]
//			|| dec_alu_transout==4'h3		//transout[15:8]
//			) ? A : 8'h00;
//	assign A_groupB = (dec_alu_input10==4'h3		//aluin10
//			|| dec_alu_input10==4'h4		//aluin11
//			|| dec_alu_input20==4'h2		//aluin20
//			|| dec_alu_input20==4'h3		//aluin21
//			|| dec_alu_mulu				//muluout
//			|| dec_alu_bitsh==5'h1c			//bitshin10
//			|| dec_alu_bitsh==5'h1d			//bitshin10
//			|| dec_alu_bitsh==5'h02			//bitshin20
//			|| dec_alu_bitsh==5'h09			//bitshin20
//			|| dec_alu_bitsh==5'h19			//bitshin20
//			|| dec_alu_bitsh==5'h0f			//bitshin20
//			|| dec_alu_bitsh==5'h03			//bitshin21
//			|| dec_movs				//Z
//			|| dec_cmps				//CY
//			) ? A : 8'h00;
//	assign A_groupC = (dec_xch_byte				//XBCDEHL��BANK0-3
//			|| dec_xchw_bc				//B��BANK0-3
//			|| dec_xchw_de				//D��BANK0-3
//			|| dec_xchw_hl				//H��BANK0-3
//			) ? A : 8'h00;
//
//	assign X_groupA = (dec_alu_transout==4'h3		//transout[7:0]
//			) ? X : 8'h00;
//	assign X_groupB = (dec_alu_transout==4'h3		//transout[7:0]
//			|| dec_alu_input10==4'h4		//aluin10
//			|| dec_alu_input20==4'h3		//aluin20
//			|| dec_alu_mulu				//muluout
//			|| dec_alu_bitsh==5'h03			//bitshin20
//			|| dec_movs				//Z
//			) ? X : 8'h00;
//	assign X_groupC = (dec_xchw_bc				//B��BANK0-3
//			|| dec_xchw_de				//D��BANK0-3
//			|| dec_xchw_hl				//H��BANK0-3
//			) ? X : 8'h00;
//
//	assign B_groupA = (dec_alu_transout==4'h4		//transout[7:0]
//			|| dec_alu_transout==4'h5		//transout[15:8]
//			) ? B : 8'h00;
//	assign B_groupB = (dec_alu_input10==4'h5		//aluin10
//			|| dec_alu_input10==4'h6		//aluin11
//			|| dec_alu_input20==4'h4		//aluin20
//			|| dec_alu_input20==4'h5		//aluin21
//			|| dec_alu_bitsh==5'h04			//bitshin20
//			|| dec_alu_bitsh==5'h05			//bitshin21
//			) ? B : 8'h00;
//	assign B_groupC = (dec_xchw_bc				//A��BANK0-3
//			) ? B : 8'h00;
//
//	assign C_groupA = (dec_alu_transout==4'h5		//transout[7:0]
//			) ? C : 8'h00;
//	assign C_groupB = (dec_alu_input10==4'h6		//aluin10
//			|| dec_alu_input20==4'h5		//aluin20
//			|| dec_alu_bitsh==5'h05			//bitshin20
//			) ? C : 8'h00;
//	assign C_groupC = (dec_xchw_bc				//X��BANK0-3
//			) ? C : 8'h00;
//
//	assign D_groupA = (dec_alu_transout==4'h6		//transout[7:0]
//			|| dec_alu_transout==4'h7		//transout[15:8]
//			) ? D : 8'h00;
//	assign D_groupB = (dec_alu_input10==4'h7		//aluin10
//			|| dec_alu_input10==4'h8		//aluin11
//			|| dec_alu_input20==4'h6		//aluin20
//			|| dec_alu_input20==4'h7		//aluin21
//			) ? D : 8'h00;
//	assign D_groupC = (dec_xchw_de				//A��BANK0-3
//			) ? D : 8'h00;
//
//	assign E_groupA = (dec_alu_transout==4'h7		//transout[7:0]
//			) ? E : 8'h00;
//	assign E_groupB = (dec_alu_input10==4'h8		//aluin10
//			|| dec_alu_input20==4'h7		//aluin20
//			) ? E : 8'h00;
//	assign E_groupC = (dec_xchw_de				//A��BANK0-3
//			) ? E : 8'h00;
//
//	assign H_groupA = (dec_alu_transout==4'h8		//transout[7:0]
//			|| dec_alu_transout==4'h9		//transout[15:8]
//			) ? H : 8'h00;
//	assign H_groupB = (dec_alu_input10==4'h9		//aluin10
//			|| dec_alu_input10==4'ha		//aluin11
//			|| dec_alu_input20==4'h8		//aluin20
//			|| dec_alu_input20==4'h9		//aluin21
//			) ? H : 8'h00;
//	assign H_groupC = (dec_xchw_hl				//A��BANK0-3
//			) ? H : 8'h00;
//
//	assign L_groupA = (dec_alu_transout==4'h9		//transout[7:0]
//			) ? L : 8'h00;
//	assign L_groupB = (dec_alu_input10==4'ha		//aluin10
//			|| dec_alu_input20==4'h9		//aluin20
//			) ? L : 8'h00;
//	assign L_groupC = (dec_xchw_hl				//A��BANK0-3
//			) ? L : 8'h00;
//
//	assign imdr_groupA = (dec_alu_transin			//transin[15:0]
//			) ? imdr : 16'h0000;
//
//	assign imdr_groupB = (dmard				//buf0, buf1
//			|| dec_alu_input10==4'hb		//aluin10, aluin11
//			|| dec_alu_input10==4'he		//aluin10, aluin11
//			|| dec_alu_input20==4'hc		//aluin20, aluin21
//			|| dec_alu_bitsh==5'h0c			//bitshin10
//			|| dec_alu_bitsh==5'h0d			//bitshin10
//			|| dec_alu_bitsh==5'h08			//bitshin20
//			|| dec_alu_bitsh==5'h18			//bitshin20
//			|| dec_alu_bitsh==5'h0e			//bitshin20
//			) ? imdr : 16'h0000;

/*------------------------------------------------------------------------------*/
// ���򤷤Ƥ���Х󥯤ȥ��ɥ쥹���ꤷ���쥸�����ΥХ󥯤����פ��Ƥ����磱�Ȥʤ롣
/*------------------------------------------------------------------------------*/
/* Ver2.0  ���ɥ쥹��vpa����ma_pre���ѹ���SLFLASH�ι�®���ΰ١�			*/
/*��������vpa�ˤ�DMA�Υ��ɥ쥹�����Ǥ��ꡢDMA�����ѥ쥸�����ؤ�ž���϶ػ�	*/
/*------------------------------------------------------------------------------*/
	assign bank_correspond = (bank0 & (ma_pre[4:3] == 2'b11)) | (bank1 & (ma_pre[4:3] == 2'b10)) |
				 (bank2 & (ma_pre[4:3] == 2'b01)) | (bank3 & (ma_pre[4:3] == 2'b00)) ;

// �ƥ쥸�����ؤΥ饤�ȥ��������ǣ��Ȥʤ롣�ϥ����ɤθ��Ф��Ѥ��롣
/*------------------------------------------------------------------------------*/
/* Ver2.0  ���ɥ쥹��vpa����ma_pre���ѹ���SLFLASH�ι�®���ΰ١�			*/
/*��������cpuwr��cpuwr_reg���ѹ���wdop��dec_word_access���ѹ���			*/
/*------------------------------------------------------------------------------*/
	assign A_access = dec_A_enable | (slreg & cpuwr_reg & bank_correspond & ((ma_pre[2:0] == 3'b001) | ({dec_word_access,ma_pre[2:0]} == 4'b1000))) ;
	assign X_access = dec_X_enable | (slreg & cpuwr_reg & bank_correspond & ( ma_pre[2:0] == 3'b000)) ;
	assign B_access = dec_B_enable | (slreg & cpuwr_reg & bank_correspond & ((ma_pre[2:0] == 3'b011) | ({dec_word_access,ma_pre[2:0]} == 4'b1010))) ;
	assign C_access = dec_C_enable | (slreg & cpuwr_reg & bank_correspond & ( ma_pre[2:0] == 3'b010)) ;
	assign D_access = dec_D_enable | (slreg & cpuwr_reg & bank_correspond & ((ma_pre[2:0] == 3'b101) | ({dec_word_access,ma_pre[2:0]} == 4'b1100))) ;
	assign E_access = dec_E_enable | (slreg & cpuwr_reg & bank_correspond & ( ma_pre[2:0] == 3'b100)) ;
	assign H_access = dec_H_enable | (slreg & cpuwr_reg & bank_correspond & ((ma_pre[2:0] == 3'b111) | ({dec_word_access,ma_pre[2:0]} == 4'b1110))) ;
	assign L_access = dec_L_enable | (slreg & cpuwr_reg & bank_correspond & ( ma_pre[2:0] == 3'b110)) ;

/*------------------------------------------------------------------------------*/
/* Ver2.0  ���ɥ쥹��vpa����ma_pre���ѹ���cpuwr��cpuwr_reg���ѹ���		*/
/*�����������ѥ쥸������_groupC���ѹ�						*/
/*------------------------------------------------------------------------------*/
// �쥸�����Х󥯣�
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) A_bank0 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait || data_hazard) A_bank0 <= A_bank0 ;
			else if (dec_A_enable & bank0) begin
				if (dec_word_access) begin
					if (dec_xchw_hl)	A_bank0 <= H_groupC ;
					else if (dec_xchw_de)	A_bank0 <= D_groupC ;
					else if (dec_xchw_bc)	A_bank0 <= B_groupC ;
					else			A_bank0 <= aluout[15:8] ;
				end
				else if (dec_xch_byte && cpuwr_reg) A_bank0 <= buf0 ;
				else				A_bank0 <= aluout[7:0] ;
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0],dec_word_access})
					({1'b1,4'h9,1'bx}) : A_bank0 <= mdw_pre[15:8] ;
					({1'b1,4'h8,1'b1}) : A_bank0 <= mdw_pre[15:8] ;
					default	: A_bank0 <= A_bank0 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) X_bank0 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait || data_hazard) X_bank0 <= X_bank0 ;
			else if (dec_X_enable & bank0) begin
				if (dec_xchw_hl)	X_bank0 <= L_groupC ;
				else if (dec_xchw_de)	X_bank0 <= E_groupC ;
				else if (dec_xchw_bc)	X_bank0 <= C_groupC ;
				else if (dec_xch_byte)	X_bank0 <= A_groupC ;
				else			X_bank0 <= aluout[7:0] ;
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0]})
					({1'b1,4'h8}) : X_bank0 <= mdw_pre[7:0] ;
					default	: X_bank0 <= X_bank0 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) B_bank0 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) B_bank0 <= B_bank0 ;
			else if (dec_B_enable & bank0) begin
				if (dec_word_access) begin
					if (dec_xchw_bc)	B_bank0 <= A_groupC ;
					else			B_bank0 <= aluout[15:8] ;
				end
				else begin
					if (dec_xch_byte)	B_bank0 <= A_groupC ;
					else			B_bank0 <= aluout[7:0] ;
				end
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0],dec_word_access})
					({1'b1,4'hb,1'bx}) : B_bank0 <= mdw_pre[15:8] ;
					({1'b1,4'ha,1'b1}) : B_bank0 <= mdw_pre[15:8] ;
					default	: B_bank0 <= B_bank0 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) C_bank0 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) C_bank0 <= C_bank0 ;
			else if (dec_C_enable & bank0) begin
				if (dec_xchw_bc)	C_bank0 <= X_groupC ;
				else if (dec_xch_byte)	C_bank0 <= A_groupC ;
				else			C_bank0 <= aluout[7:0] ;
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0]})
					({1'b1,4'ha}) : C_bank0 <= mdw_pre[7:0] ;
					default	: C_bank0 <= C_bank0 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) D_bank0 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) D_bank0 <= D_bank0 ;
			else if (dec_D_enable & bank0) begin
				if (dec_word_access) begin
					if (dec_xchw_de)	D_bank0 <= A_groupC ;
					else			D_bank0 <= aluout[15:8] ;
				end
				else begin
					if (dec_xch_byte)	D_bank0 <= A_groupC ;
					else			D_bank0 <= aluout[7:0] ;
				end
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0],dec_word_access})
					({1'b1,4'hd,1'bx}) : D_bank0 <= mdw_pre[15:8] ;
					({1'b1,4'hc,1'b1}) : D_bank0 <= mdw_pre[15:8] ;
					default	: D_bank0 <= D_bank0 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) E_bank0 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) E_bank0 <= E_bank0 ;
			else if (dec_E_enable & bank0) begin
				if (dec_xchw_de)	E_bank0 <= X_groupC ;
				else if (dec_xch_byte)	E_bank0 <= A_groupC ;
				else			E_bank0 <= aluout[7:0] ;
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0]})
					({1'b1,4'hc}) : E_bank0 <= mdw_pre[7:0] ;
					default	: E_bank0 <= E_bank0 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) H_bank0 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) H_bank0 <= H_bank0 ;
			else if (dec_H_enable & bank0) begin
				if (dec_word_access) begin
					if (dec_xchw_hl)	H_bank0 <= A_groupC ;
					else			H_bank0 <= aluout[15:8] ;
				end
				else begin
					if (dec_xch_byte)	H_bank0 <= A_groupC ;
					else			H_bank0 <= aluout[7:0] ;
				end
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0],dec_word_access})
					({1'b1,4'hf,1'bx}) : H_bank0 <= mdw_pre[15:8] ;
					({1'b1,4'he,1'b1}) : H_bank0 <= mdw_pre[15:8] ;
					default	: H_bank0 <= H_bank0 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) L_bank0 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) L_bank0 <= L_bank0 ;
			else if (dec_L_enable & bank0) begin
				if (dec_xchw_hl)	L_bank0 <= X_groupC ;
				else if (dec_xch_byte)	L_bank0 <= A_groupC ;
				else			L_bank0 <= aluout[7:0] ;
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0]})
					({1'b1,4'he}) : L_bank0 <= mdw_pre[7:0] ;
					default	: L_bank0 <= L_bank0 ;
				endcase
			end
		end
	end

// �쥸�����Х󥯣�
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) A_bank1 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait || data_hazard) A_bank1 <= A_bank1 ;
			else if (dec_A_enable & bank1) begin
				if (dec_word_access) begin
					if (dec_xchw_hl)	A_bank1 <= H_groupC ;
					else if (dec_xchw_de)	A_bank1 <= D_groupC ;
					else if (dec_xchw_bc)	A_bank1 <= B_groupC ;
					else			A_bank1 <= aluout[15:8] ;
				end
				else if (dec_xch_byte && cpuwr_reg) A_bank1 <= buf0 ;
				else				A_bank1 <= aluout[7:0] ;
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0],dec_word_access})
					({1'b1,4'h1,1'bx}) : A_bank1 <= mdw_pre[15:8] ;
					({1'b1,4'h0,1'b1}) : A_bank1 <= mdw_pre[15:8] ;
					default	: A_bank1 <= A_bank1 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) X_bank1 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait || data_hazard) X_bank1 <= X_bank1 ;
			else if (dec_X_enable & bank1) begin
				if (dec_xchw_hl)	X_bank1 <= L_groupC ;
				else if (dec_xchw_de)	X_bank1 <= E_groupC ;
				else if (dec_xchw_bc)	X_bank1 <= C_groupC ;
				else if (dec_xch_byte)	X_bank1 <= A_groupC ;
				else			X_bank1 <= aluout[7:0] ;
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0]})
					({1'b1,4'h0}) : X_bank1 <= mdw_pre[7:0] ;
					default	: X_bank1 <= X_bank1 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) B_bank1 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) B_bank1 <= B_bank1 ;
			else if (dec_B_enable & bank1) begin
				if (dec_word_access) begin
					if (dec_xchw_bc)	B_bank1 <= A_groupC ;
					else			B_bank1 <= aluout[15:8] ;
				end
				else begin
					if (dec_xch_byte)	B_bank1 <= A_groupC ;
					else			B_bank1 <= aluout[7:0] ;
				end
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0],dec_word_access})
					({1'b1,4'h3,1'bx}) : B_bank1 <= mdw_pre[15:8] ;
					({1'b1,4'h2,1'b1}) : B_bank1 <= mdw_pre[15:8] ;
					default	: B_bank1 <= B_bank1 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) C_bank1 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) C_bank1 <= C_bank1 ;
			else if (dec_C_enable & bank1) begin
				if (dec_xchw_bc)	C_bank1 <= X_groupC ;
				else if (dec_xch_byte)	C_bank1 <= A_groupC ;
				else			C_bank1 <= aluout[7:0] ;
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0]})
					({1'b1,4'h2}) : C_bank1 <= mdw_pre[7:0] ;
					default	: C_bank1 <= C_bank1 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) D_bank1 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) D_bank1 <= D_bank1 ;
			else if (dec_D_enable & bank1) begin
				if (dec_word_access) begin
					if (dec_xchw_de)	D_bank1 <= A_groupC ;
					else			D_bank1 <= aluout[15:8] ;
				end
				else begin
					if (dec_xch_byte)	D_bank1 <= A_groupC ;
					else			D_bank1 <= aluout[7:0] ;
				end
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0],dec_word_access})
					({1'b1,4'h5,1'bx}) : D_bank1 <= mdw_pre[15:8] ;
					({1'b1,4'h4,1'b1}) : D_bank1 <= mdw_pre[15:8] ;
					default	: D_bank1 <= D_bank1 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) E_bank1 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) E_bank1 <= E_bank1 ;
			else if (dec_E_enable & bank1) begin
				if (dec_xchw_de)	E_bank1 <= X_groupC ;
				else if (dec_xch_byte)	E_bank1 <= A_groupC ;
				else			E_bank1 <= aluout[7:0] ;
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0]})
					({1'b1,4'h4}) : E_bank1 <= mdw_pre[7:0] ;
					default	: E_bank1 <= E_bank1 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) H_bank1 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) H_bank1 <= H_bank1 ;
			else if (dec_H_enable & bank1) begin
				if (dec_word_access) begin
					if (dec_xchw_hl)	H_bank1 <= A_groupC ;
					else			H_bank1 <= aluout[15:8] ;
				end
				else begin
					if (dec_xch_byte)	H_bank1 <= A_groupC ;
					else			H_bank1 <= aluout[7:0] ;
				end
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0],dec_word_access})
					({1'b1,4'h7,1'bx}) : H_bank1 <= mdw_pre[15:8] ;
					({1'b1,4'h6,1'b1}) : H_bank1 <= mdw_pre[15:8] ;
					default	: H_bank1 <= H_bank1 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) L_bank1 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) L_bank1 <= L_bank1 ;
			else if (dec_L_enable & bank1) begin
				if (dec_xchw_hl)	L_bank1 <= X_groupC ;
				else if (dec_xch_byte)	L_bank1 <= A_groupC ;
				else			L_bank1 <= aluout[7:0] ;
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0]})
					({1'b1,4'h6}) : L_bank1 <= mdw_pre[7:0] ;
					default	: L_bank1 <= L_bank1 ;
				endcase
			end
		end
	end

// �쥸�����Х󥯣�
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) A_bank2 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait || data_hazard) A_bank2 <= A_bank2 ;
			else if (dec_A_enable & bank2) begin
				if (dec_word_access) begin
					if (dec_xchw_hl)	A_bank2 <= H_groupC ;
					else if (dec_xchw_de)	A_bank2 <= D_groupC ;
					else if (dec_xchw_bc)	A_bank2 <= B_groupC ;
					else			A_bank2 <= aluout[15:8] ;
				end
				else if (dec_xch_byte && cpuwr_reg) A_bank2 <= buf0 ;
				else				A_bank2 <= aluout[7:0] ;
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0],dec_word_access})
					({1'b0,4'h9,1'bx}) : A_bank2 <= mdw_pre[15:8] ;
					({1'b0,4'h8,1'b1}) : A_bank2 <= mdw_pre[15:8] ;
					default	: A_bank2 <= A_bank2 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) X_bank2 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait || data_hazard) X_bank2 <= X_bank2 ;
			else if (dec_X_enable & bank2) begin
				if (dec_xchw_hl)	X_bank2 <= L_groupC ;
				else if (dec_xchw_de)	X_bank2 <= E_groupC ;
				else if (dec_xchw_bc)	X_bank2 <= C_groupC ;
				else if (dec_xch_byte)	X_bank2 <= A_groupC ;
				else			X_bank2 <= aluout[7:0] ;
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0]})
					({1'b0,4'h8}) : X_bank2 <= mdw_pre[7:0] ;
					default	: X_bank2 <= X_bank2 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) B_bank2 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) B_bank2 <= B_bank2 ;
			else if (dec_B_enable & bank2) begin
				if (dec_word_access) begin
					if (dec_xchw_bc)	B_bank2 <= A_groupC ;
					else			B_bank2 <= aluout[15:8] ;
				end
				else begin
					if (dec_xch_byte)	B_bank2 <= A_groupC ;
					else			B_bank2 <= aluout[7:0] ;
				end
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0],dec_word_access})
					({1'b0,4'hb,1'bx}) : B_bank2 <= mdw_pre[15:8] ;
					({1'b0,4'ha,1'b1}) : B_bank2 <= mdw_pre[15:8] ;
					default	: B_bank2 <= B_bank2 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) C_bank2 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) C_bank2 <= C_bank2 ;
			else if (dec_C_enable & bank2) begin
				if (dec_xchw_bc)	C_bank2 <= X_groupC ;
				else if (dec_xch_byte)	C_bank2 <= A_groupC ;
				else			C_bank2 <= aluout[7:0] ;
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0]})
					({1'b0,4'ha}) : C_bank2 <= mdw_pre[7:0] ;
					default	: C_bank2 <= C_bank2 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) D_bank2 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) D_bank2 <= D_bank2 ;
			else if (dec_D_enable & bank2) begin
				if (dec_word_access) begin
					if (dec_xchw_de)	D_bank2 <= A_groupC ;
					else			D_bank2 <= aluout[15:8] ;
				end
				else begin
					if (dec_xch_byte)	D_bank2 <= A_groupC ;
					else			D_bank2 <= aluout[7:0] ;
				end
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0],dec_word_access})
					({1'b0,4'hd,1'bx}) : D_bank2 <= mdw_pre[15:8] ;
					({1'b0,4'hc,1'b1}) : D_bank2 <= mdw_pre[15:8] ;
					default	: D_bank2 <= D_bank2 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) E_bank2 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) E_bank2 <= E_bank2 ;
			else if (dec_E_enable & bank2) begin
				if (dec_xchw_de)	E_bank2 <= X_groupC ;
				else if (dec_xch_byte)	E_bank2 <= A_groupC ;
				else			E_bank2 <= aluout[7:0] ;
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0]})
					({1'b0,4'hc}) : E_bank2 <= mdw_pre[7:0] ;
					default	: E_bank2 <= E_bank2 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) H_bank2 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) H_bank2 <= H_bank2 ;
			else if (dec_H_enable & bank2) begin
				if (dec_word_access) begin
					if (dec_xchw_hl)	H_bank2 <= A_groupC ;
					else			H_bank2 <= aluout[15:8] ;
				end
				else begin
					if (dec_xch_byte)	H_bank2 <= A_groupC ;
					else			H_bank2 <= aluout[7:0] ;
				end
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0],dec_word_access})
					({1'b0,4'hf,1'bx}) : H_bank2 <= mdw_pre[15:8] ;
					({1'b0,4'he,1'b1}) : H_bank2 <= mdw_pre[15:8] ;
					default	: H_bank2 <= H_bank2 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) L_bank2 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) L_bank2 <= L_bank2 ;
			else if (dec_L_enable & bank2) begin
				if (dec_xchw_hl)	L_bank2 <= X_groupC ;
				else if (dec_xch_byte)	L_bank2 <= A_groupC ;
				else			L_bank2 <= aluout[7:0] ;
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0]})
					({1'b0,4'he}) : L_bank2 <= mdw_pre[7:0] ;
					default	: L_bank2 <= L_bank2 ;
				endcase
			end
		end
	end

// �쥸�����Х󥯣�
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) A_bank3 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait || data_hazard) A_bank3 <= A_bank3 ;
			else if (dec_A_enable & bank3) begin
				if (dec_word_access) begin
					if (dec_xchw_hl)	A_bank3 <= H_groupC ;
					else if (dec_xchw_de)	A_bank3 <= D_groupC ;
					else if (dec_xchw_bc)	A_bank3 <= B_groupC ;
					else			A_bank3 <= aluout[15:8] ;
				end
				else if (dec_xch_byte && cpuwr_reg) A_bank3 <= buf0 ;
				else				A_bank3 <= aluout[7:0] ;
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0],dec_word_access})
					({1'b0,4'h1,1'bx}) : A_bank3 <= mdw_pre[15:8] ;
					({1'b0,4'h0,1'b1}) : A_bank3 <= mdw_pre[15:8] ;
					default	: A_bank3 <= A_bank3 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) X_bank3 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait || data_hazard) X_bank3 <= X_bank3 ;
			else if (dec_X_enable & bank3) begin
				if (dec_xchw_hl)	X_bank3 <= L_groupC ;
				else if (dec_xchw_de)	X_bank3 <= E_groupC ;
				else if (dec_xchw_bc)	X_bank3 <= C_groupC ;
				else if (dec_xch_byte)	X_bank3 <= A_groupC ;
				else			X_bank3 <= aluout[7:0] ;
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0]})
					({1'b0,4'h0}) : X_bank3 <= mdw_pre[7:0] ;
					default	: X_bank3 <= X_bank3 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) B_bank3 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) B_bank3 <= B_bank3 ;
			else if (dec_B_enable & bank3) begin
				if (dec_word_access) begin
					if (dec_xchw_bc)	B_bank3 <= A_groupC ;
					else			B_bank3 <= aluout[15:8] ;
				end
				else begin
					if (dec_xch_byte)	B_bank3 <= A_groupC ;
					else			B_bank3 <= aluout[7:0] ;
				end
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0],dec_word_access})
					({1'b0,4'h3,1'bx}) : B_bank3 <= mdw_pre[15:8] ;
					({1'b0,4'h2,1'b1}) : B_bank3 <= mdw_pre[15:8] ;
					default	: B_bank3 <= B_bank3 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) C_bank3 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) C_bank3 <= C_bank3 ;
			else if (dec_C_enable & bank3) begin
				if (dec_xchw_bc)	C_bank3 <= X_groupC ;
				else if (dec_xch_byte)	C_bank3 <= A_groupC ;
				else			C_bank3 <= aluout[7:0] ;
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0]})
					({1'b0,4'h2}) : C_bank3 <= mdw_pre[7:0] ;
					default	: C_bank3 <= C_bank3 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) D_bank3 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) D_bank3 <= D_bank3 ;
			else if (dec_D_enable & bank3) begin
				if (dec_word_access) begin
					if (dec_xchw_de)	D_bank3 <= A_groupC ;
					else			D_bank3 <= aluout[15:8] ;
				end
				else begin
					if (dec_xch_byte)	D_bank3 <= A_groupC ;
					else			D_bank3 <= aluout[7:0] ;
				end
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0],dec_word_access})
					({1'b0,4'h5,1'bx}) : D_bank3 <= mdw_pre[15:8] ;
					({1'b0,4'h4,1'b1}) : D_bank3 <= mdw_pre[15:8] ;
					default	: D_bank3 <= D_bank3 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) E_bank3 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) E_bank3 <= E_bank3 ;
			else if (dec_E_enable & bank3) begin
				if (dec_xchw_de)	E_bank3 <= X_groupC ;
				else if (dec_xch_byte)	E_bank3 <= A_groupC ;
				else			E_bank3 <= aluout[7:0] ;
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0]})
					({1'b0,4'h4}) : E_bank3 <= mdw_pre[7:0] ;
					default	: E_bank3 <= E_bank3 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) H_bank3 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) H_bank3 <= H_bank3 ;
			else if (dec_H_enable & bank3) begin
				if (dec_word_access) begin
					if (dec_xchw_hl)	H_bank3 <= A_groupC ;
					else			H_bank3 <= aluout[15:8] ;
				end
				else begin
					if (dec_xch_byte)	H_bank3 <= A_groupC ;
					else			H_bank3 <= aluout[7:0] ;
				end
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0],dec_word_access})
					({1'b0,4'h7,1'bx}) : H_bank3 <= mdw_pre[15:8] ;
					({1'b0,4'h6,1'b1}) : H_bank3 <= mdw_pre[15:8] ;
					default	: H_bank3 <= H_bank3 ;
				endcase
			end
		end
	end

	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) L_bank3 <= 8'h00 ;
// for EVA
//		else if (cpuen) begin
                else if (cpuen & ~sel_svmod_reg) begin
//
			if (reg_wait) L_bank3 <= L_bank3 ;
			else if (dec_L_enable & bank3) begin
				if (dec_xchw_hl)	L_bank3 <= X_groupC ;
				else if (dec_xch_byte)	L_bank3 <= A_groupC ;
				else			L_bank3 <= aluout[7:0] ;
			end
			else if (slreg && cpuwr_reg) begin
				casex ({ma_pre[4:0]})
					({1'b0,4'h6}) : L_bank3 <= mdw_pre[7:0] ;
					default	: L_bank3 <= L_bank3 ;
				endcase
			end
		end
	end

// for EVA
// for SVMODE

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb) A_sv <= 8'h00 ;
                else if (cpuen & sel_svmod_reg) begin
                        if (reg_wait || data_hazard) A_sv <= A ;
                        else if (dec_A_enable) begin
                                if (dec_word_access) begin
                                        if (dec_xchw_hl)        A_sv <= H ;
                                        else if (dec_xchw_de)   A_sv <= D ;
                                        else if (dec_xchw_bc)   A_sv <= B ;
                                        else                    A_sv <= aluout[15:8] ;
                                end
                                else if (dec_xch_byte && cpuwr) A_sv <= buf0 ;
                                else                            A_sv <= aluout[7:0] ;
                        end
                end
        end

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb) X_sv <= 8'h00 ;
                else if (cpuen & sel_svmod_reg) begin
                        if (reg_wait || data_hazard) X_sv <= X ;
                        else if (dec_X_enable) begin
                                if (dec_xchw_hl)        X_sv <= L ;
                                else if (dec_xchw_de)   X_sv <= E ;
                                else if (dec_xchw_bc)   X_sv <= C ;
                                else if (dec_xch_byte)  X_sv <= A ;
                                else                    X_sv <= aluout[7:0] ;
                        end     
                end
        end

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb) B_sv <= 8'h00 ;
                else if (cpuen & sel_svmod_reg) begin
                        if (reg_wait) B_sv <= B ;
                        else if (dec_B_enable) begin
                                if (dec_word_access) begin
                                        if (dec_xchw_bc)        B_sv <= A ;
                                        else                    B_sv <= aluout[15:8] ;
                                end
                                else begin
                                        if (dec_xch_byte)       B_sv <= A ;
                                        else                    B_sv <= aluout[7:0] ;
                                end
                        end
                end
        end

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb) C_sv <= 8'h00 ;
                else if (cpuen & sel_svmod_reg) begin
                        if (reg_wait) C_sv <= C ;
                        else if (dec_C_enable) begin
                                if (dec_xchw_bc)        C_sv <= X ;
                                else if (dec_xch_byte)  C_sv <= A ;
                                else                    C_sv <= aluout[7:0] ;
                        end
                end
        end

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb) D_sv <= 8'h00 ;
                else if (cpuen & sel_svmod_reg) begin
                        if (reg_wait) D_sv <= D ;
                        else if (dec_D_enable) begin
                                if (dec_word_access) begin
                                        if (dec_xchw_de)        D_sv <= A ;
                                        else                    D_sv <= aluout[15:8] ;
                                end
                                else begin
                                        if (dec_xch_byte)       D_sv <= A ;
                                        else                    D_sv <= aluout[7:0] ;
                                end
                        end
                end
        end

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb) E_sv <= 8'h00 ;
                else if (cpuen & sel_svmod_reg) begin
                        if (reg_wait) E_sv <= E ;
                        else if (dec_E_enable) begin
                                if (dec_xchw_de)        E_sv <= X ;
                                else if (dec_xch_byte)  E_sv <= A ;
                                else                    E_sv <= aluout[7:0] ;
                        end
                end
        end

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb) H_sv <= 8'h00 ;
                else if (cpuen & sel_svmod_reg) begin
                        if (reg_wait) H_sv <= H ;
                        else if (dec_H_enable) begin
                                if (dec_word_access) begin
                                        if (dec_xchw_hl)        H_sv <= A ;
                                        else                    H_sv <= aluout[15:8] ;
                                end
                                else begin
                                        if (dec_xch_byte)       H_sv <= A ;
                                        else                    H_sv <= aluout[7:0] ;
                                end
                        end
                end
        end

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb) L_sv <= 8'h00 ;
                else if (cpuen & sel_svmod_reg) begin
                        if (reg_wait) L_sv <= L ;
                        else if (dec_L_enable) begin
                                if (dec_xchw_hl)        L_sv <= X ;
                                else if (dec_xch_byte)  L_sv <= A ;
                                else                    L_sv <= aluout[7:0] ;
                        end
                end
        end
//

/*------------------------------------------------------------------------------*/
/* �ǡ����ݻ��Хåե�								*/
/*------------------------------------------------------------------------------*/
/*   �أã�̿�ᡢ�����å�ư�������ȯ�������˥ǡ������ݻ����롣		*/
/*------------------------------------------------------------------------------*/

// ma�β��̣��ӥå�maw1���ɤ߽Ф�PID�Υǡ��������򤹤롣
/*------------------------------------------------------------------------------*/
/* Ver2.0  Flash�ɤ߽Ф����Ƥ��ʤ�����rdata�򣰤˸��ꡣ				*/
/*------------------------------------------------------------------------------*/
	always @(maw1 or pid or pa_data_buf) begin
		if (maw1)	rdata = pid[31:16] ;
		else		rdata = pid[15:0] ;
//		if (pa_data_buf) begin
//			if (maw1)	rdata = pid[31:16] ;
//			else		rdata = pid[15:0] ;
//		end
//		else rdata = 8'h00;
	end

// �ǡ����ݻ��Хåե����̣��ӥå�
// XCH̿�ᡢ�����å�ư�������ȯ������FLASH�꡼�ɥ�����������DMAž������
// buf0�쥸����������ǡ��������򤹤롣
/*------------------------------------------------------------------------------*/
/* Ver2.0  bufr��ɬ�פʻ���������_groupB���ѹ�					*/
/*------------------------------------------------------------------------------*/
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) buf0 <= 8'h00 ;
		else if (cpuen || waitdma) begin
			if (dmard && vpa[0])			buf0 <= imdr_groupB[15:8] ;
			else if (dmard && !vpa[0])		buf0 <= imdr_groupB[7:0] ;
			else if (reg_wait && !pa_data_buf)	buf0 <= buf0 ;
			else if (dec_buf0_enable || dmard || dec_set_buf_retadr || dec_set_buf_intr || pa_data_buf) begin
				if (dec_set_buf_retadr)		buf0 <= pc_inc[7:0] ;
				else if (dec_set_buf_intr)	buf0 <= pc[7:0] ;
				else if (pa_data_buf)		buf0 <= rdata[7:0] ;
				else				buf0 <= aluout[7:0] ;
			end
		end
	end

// �ǡ����ݻ��Хåե���̣��ӥå�
// XCH̿�ᡢ�����å�ư�������ȯ������FLASH�꡼�ɥ�����������DMAž������
// buf1�쥸����������ǡ��������򤹤롣
/*------------------------------------------------------------------------------*/
/* Ver2.0  bufr��ɬ�פʻ���������_groupB���ѹ�					*/
/*------------------------------------------------------------------------------*/
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) buf1 <= 8'h00 ;
		else if (cpuen || waitdma) begin
			if (dmard && vpa[0])			buf1 <= imdr_groupB[7:0] ;
			else if (dmard && !vpa[0])		buf1 <= imdr_groupB[15:8] ;
			else if (reg_wait && !pa_data_buf)	buf1 <= buf1 ;
			else if (dec_buf1_enable || dmard || dec_set_buf_retadr || dec_set_buf_intr || pa_data_buf) begin
				if (dec_set_buf_retadr)		buf1 <= pc_inc[15:8] ;
				else if (dec_set_buf_intr)	buf1 <= pc[15:8] ;
				else if (pa_data_buf)		buf1 <= rdata[15:8] ;
				else				buf1 <= aluout[15:8] ;
			end
		end
	end

// ���������ݻ��Хåե�
// XCH̿�ᡢ�����å�ư�������ȯ������buf2�쥸����������ǡ��������򤹤롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) buf2 <= 4'h0 ;
		else if (cpuen) begin
			if (reg_wait) buf2 <= buf2 ;
			else if (dec_buf2_enable || dec_set_buf_retadr || dec_set_buf_intr) begin
				if (dec_set_buf_retadr)		buf2 <= pc_inc[19:16] ;
				else if (dec_set_buf_intr)	buf2 <= pc[19:16] ;
				else				buf2 <= aluout[3:0] ;
			end
		end
	end

/*------------------------------------------------------------------------------*/
/* �����å��ݥ���								*/
/*------------------------------------------------------------------------------*/
/*   �����å����줿�ǡ����Υ��ɥ쥹�򼨤���					*/
/*------------------------------------------------------------------------------*/

// �ǥ�������������濮��ˤ��SP��ǥ�����Ȥ��뤫���󥯥���Ȥ��뤫������
	always @(SP or dec_sp_dec or dec_sp_inc) begin
		if (dec_sp_dec)		sp_pre = SP + 15'h7fff ;
		else if (dec_sp_inc)	sp_pre = SP + 15'h0001 ;
		else			sp_pre = SP ;
	end

// �����å�ư����Υ��ꥢ�ɥ쥹��
// ������ȯ���������ߤ�SP�ͤȥǥ�����ȸ��SP�ͤ���ꥢ�ɥ쥹�Ȥ��ƽ��Ϥ��롣
	assign sp_inc = (dec_sp_dec) ? sp_pre : SP ;

// for EVA

        reg             spinc, spdec;

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb) begin
                        spinc <= 1'b0 ;
                        spdec <= 1'b0 ;
                        end
                else if (cpuen) begin
                        if (reg_wait) begin
                                spinc <= spinc ;
                                spdec <= spdec ;
                        end
                        else if (data_hazard_flg) begin
                                spinc <= spinc ;
                                spdec <= spdec ;
                        end
                        else begin
                                spinc <= dec_sp_inc ;
                                spdec <= dec_sp_dec ;
                        end
                end
        end
//

// �����å��ݥ��󥿡�FLASH�ե��å��ʳ��������������Ȥ�ȯ����������
// RAM�ե��å��ʳ��ǥϥ����ɰʳ��������������Ȥ�ȯ��������硢
// ������������ȯ�����ʳ���̿��μ¹Ծ��֤˰ܹԤ������RAM�ե��å����FLASH���֤򥢥�������������ݻ�����롣
// �����ؤ���ȡ������å�ư����˥������Ȥ�ȯ����������SP�����Ѥ�äƤϤ����ʤ���
// ��������FLASH�Υǡ�����������ľ���ʬ��������ϡ��㳰�Ȥ���SP�����Ѥ����������
// reg_wait�ˤ�륦�����Ȥϴ���Ū�ˤ�FLASH�ե��å����̵���Ȥʤ뤬��SP�񤭴����ȶ��礷�����ϡ�ͭ���ˤ��롣
// ID���ơ������ݻ���郎��MEM���ơ����ι�����˸���Ƥʤ��ͤ�pc_wait_flg�˴ط�������ϡ�SP������������ǥޥ������롣
// for EVA
////	//synopsys async_set_reset "resb"
////	always @(posedge baseck or negedge resb) begin
////		if (!resb)					SP <= 15'h7e00 ;
////		else if (cpuen) begin
////			if ((reg_wait && !((slflash & ~SP_enable) || pa_data_spen || sp_hazard)) ||
////			    (((!fchiram && (!data_hazard_flg && pc_wait_flg)) || (pa_st2 && !pc_wait_flg) ||
////			     (fchiram && (slflash || (slmirr && dec_sp_inc)) && pc_wait_flg)) && !SP_enable))	SP <= SP ;
////			else if (dec_SP_enable)						SP <= aluout[15:1] ;
////			else if (pselcpu && cpuwr && (vpa[3:1] == 3'b100)) begin
////				casex ({vpa[0],wdop})
////					({1'b0,1'b0}) : SP <= {SP[14:7],mdw_pre[7:1]} ;
////					({1'b0,1'b1}) : SP <= mdw_pre[15:1] ;
////					({1'b1,1'bx}) : SP <= {mdw_pre[15:8],SP[6:0]} ;
////					// cannot reach DEFAULT brunch
////					// default	: SP <= SP ;
////				endcase
////			end
////			else if (dec_sp_set_enable && (!data_hazard_flg || fchiram))	SP <= sp_pre ;
////		end
////	end
// for EVA

        assign SP0 = 1'b0 ;

        output  [14:0]  SP_usr, SP_sv;
        reg     [14:0]  SP_usr, SP_sv;

        wire svmod_sp = (svmod | svmodi) & ~(alt1) ;

        assign SP = (svmod_sp) ? SP_sv : SP_usr ;

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb)                                      SP_usr <= 15'h7e00 ;
                else if (cpuen & ~svmod_sp) begin
                        if ((reg_wait && !((slflash & !SP_enable) || pa_data_spen || sp_hazard)) ||
                            (((!fchiram && (!data_hazard_flg && pc_wait_flg)) || (pa_st2 && !pc_wait_flg) ||
                             (fchiram && (slflash || (slmirr && dec_sp_inc)) && pc_wait_flg)) && !SP_enable))   SP_usr <= SP ;
                        else if (dec_SP_enable)                                         SP_usr <= aluout[15:1] ;
                        else if (pselcpu && cpuwr && (vpa[3:1] == 3'b100)) begin
                                casex ({vpa[0],wdop})
                                        ({1'b0,1'b0}) : SP_usr <= {SP[14:7],mdw_pre[7:1]} ;
                                        ({1'b0,1'b1}) : SP_usr <= mdw_pre[15:1] ;
                                        ({1'b1,1'bx}) : SP_usr <= {mdw_pre[15:8],SP[6:0]} ;
                                // cannot reach DEFAULT brunch
                                // default      : SP_usr <= SP ;
                                endcase
                        end
                        else if (dec_sp_set_enable && (!data_hazard_flg || fchiram))    SP_usr <= sp_pre ;
                end
        end

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb)                                      SP_sv <= 15'h7f00 ;
                else if (cpuen & svmod_sp) begin
                        if ((reg_wait && !((slflash & !SP_enable) || pa_data_spen || sp_hazard)) ||
                            (((!fchiram && (!data_hazard_flg && pc_wait_flg)) || (pa_st2 && !pc_wait_flg) ||
                             (fchiram && (slflash || (slmirr && dec_sp_inc)) && pc_wait_flg)) && !SP_enable))   SP_sv <= SP ;
                        else if (dec_SP_enable)                                         SP_sv <= aluout[15:1] ;
                        else if (pselcpu && cpuwr && (vpa[3:1] == 3'b100)) begin
                                casex ({vpa[0],wdop})
                                        ({1'b0,1'b0}) : SP_sv <= {SP[14:7],mdw_pre[7:1]} ;
                                        ({1'b0,1'b1}) : SP_sv <= mdw_pre[15:1] ;
                                        ({1'b1,1'bx}) : SP_sv <= {mdw_pre[15:8],SP[6:0]} ;
                                        // cannot reach DEFAULT brunch
                                        // default      : SP_sv <= SP ;
                                endcase
                        end
                        else if (dec_sp_set_enable && (!data_hazard_flg || fchiram))    SP_sv <= sp_pre ;
                end
        end
//

// SP�ؤΥ���������ɽ�����档
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) sp_sfr_msk <= 1'b0 ;
		else if (cpuen) begin
			if (reg_wait) begin
				sp_sfr_msk <= sp_sfr_msk ;
			end
			else begin
				sp_sfr_msk <= dec_sp_set_enable & ((sp_inc[14:7] == 8'hff) | (sp_inc[14:10] == {4'h0,1'b0}) |
								   (sp_inc[14:9] == {4'h0,2'b10}) |
								   ({sp_inc[14:7],sp_inc[6:4]} == {8'hfe,3'h7})) ;
			end
		end
	end

// SP�˥����������륿���ߥ󥰤ǡ�SP��SFR���֤�ؤ�����磱�Ȥʤ롣
	assign sp_sfr_en = sp_sfr_msk ;

/*------------------------------------------------------------------------------*/
/* ����ؤΥ饤�ȥǡ���							*/
/*------------------------------------------------------------------------------*/
/*   �ǡ�������ؤΥ饤�ȥǡ������������롣					*/
/*------------------------------------------------------------------------------*/

// ��ɥ����������档��ɥ����������������RAM�ե��å���ϣ���
// RAM�ե��å����RAM�ǡ�������������ȯ����������Ω�������롣
// DMAž������dmawdop�����򤵤�롣
	assign wdop_pre = dec_word_access | (~(cpuwr | fchiram_cpurd | pa_data_mem) & fchiram) ;
	assign wdop = (waitdma) ? dmawdop : wdop_pre ;

// ��ɥǡ����Υ饤�ȥ��������ǣ��Ȥʤ롣RAM�����������ѿ��档
	assign wdwr = wdop & cpuwr ;

// ����饤�ȥǡ�������ɥ��������ξ���ALU���ϡ�
// �Х��ȥ��������ξ��ϥ��ꥢ�ɥ쥹�κǲ��̥ӥåȤ�ALU���Ϥ�ɤ���˽Ф������򤹤롣
// DMAž����ϥǡ����ݻ��Хåե������򤵤�롣
/*------------------------------------------------------------------------------*/
/* Ver2.0  MDW�ؤν��Ϥ����Ѥǿ��ߤ���transout����Ϥ��롣			*/
/*------------------------------------------------------------------------------*/
	assign mdw_pre = (wdop_pre) ? transout : (vpa[0]) ? {transout[7:0],8'h00} : {8'h00,transout[7:0]} ;
	assign mdw_dma = (dmawdop) ? {buf1,buf0} : (vpa[0]) ? {buf0,8'h00} : {8'h00,buf0} ;

	assign mdw = (dmawr) ? mdw_dma : mdw_pre ;

/*------------------------------------------------------------------------------*/
/* ��ĥ�ǡ����������ȥ쥸���� �ţ�						*/
/*------------------------------------------------------------------------------*/
/*   ̿�����إ꡼�ɥ������������Ѥ��롣					*/
/*------------------------------------------------------------------------------*/

// ���ꥢ�ɥ쥹���ղä���FLASH�������˥ǡ������������Ǥ���褦�ˤ��롣
// for EVA
////	//synopsys async_set_reset "resb"
////	always @(posedge baseck or negedge resb) begin
////		if (!resb)		ES <= 4'hf ;
////		else if (cpuen) begin
////			if (reg_wait)	ES <= ES ;
////			else if (dec_ES_enable)	ES <= aluout[3:0] ;
////			else if (pselcpu && cpuwr) begin
////				casex ({vpa,wdop})
////					({4'hc,1'b1}) : ES <= mdw_pre[11:8] ;
////					({4'hd,1'bx}) : ES <= mdw_pre[11:8] ;
////					default	: ES <= ES ;
////				endcase
////			end
////		end
////	end
// for EVA

        reg     [3:0]   ES_usr, ES_sv;

        assign ES = (sel_svmod_reg) ? ES_sv : ES_usr ;

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb)              ES_usr <= 4'hf ;
                else if (cpuen && !sel_svmod_reg) begin
                        if (reg_wait)   ES_usr <= ES ;
                        else if (dec_ES_enable) ES_usr <= aluout[3:0] ;
                        else if (pselcpu && cpuwr) begin
                                casex ({vpa,wdop})
                                        ({4'hc,1'b1}) : ES_usr <= mdw_pre[11:8] ;
                                        ({4'hd,1'bx}) : ES_usr <= mdw_pre[11:8] ;
                                        default : ES_usr <= ES ;
                                endcase
                        end
                end
        end

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb)              ES_sv <= 4'hf ;
                else if (cpuen && sel_svmod_reg) begin
                        if (reg_wait)   ES_sv <= ES ;
                        else if (dec_ES_enable) ES_sv <= aluout[3:0] ;
                        else if (pselcpu && cpuwr) begin
                                casex ({vpa,wdop})
                                        ({4'hc,1'b1}) : ES_sv <= mdw_pre[11:8] ;
                                        ({4'hd,1'bx}) : ES_sv <= mdw_pre[11:8] ;
                                        default : ES_sv <= ES ;
                                endcase
                        end
                end
        end
//

/*------------------------------------------------------------------------------*/
/* �����ɥ������ȥ쥸���� �ã�						*/
/*------------------------------------------------------------------------------*/
/*   �ǡ�������ؤΥե��å��������������Ѥ��롣				*/
/*------------------------------------------------------------------------------*/
/* Ver2.0  CS�ؤν񤭹��ߤ�CS_enable����Ѥ��ƽ񤭹���				*/
/*------------------------------------------------------------------------------*/

// �ץ���ॢ�ɥ쥹���ղä���RAM���֤˥ե��å����������Ǥ����ͤˤʤ롣
// for EVA
////	//synopsys async_set_reset "resb"
////	always @(posedge baseck or negedge resb) begin
////		if (!resb)		CS <= 4'h0 ;
////		else if (cpuen) begin
////			if (reg_wait)	CS <= CS ;
////			else if (CS_enable) CS <= mdw_pre[3:0] ;
////		end
////	end
// for EVA

        reg     [3:0]   CS_usr, CS_sv;

        assign CS = (sel_svmod_reg) ? CS_sv : CS_usr ;

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb)              CS_usr <= 4'h0 ;
                else if (cpuen && !sel_svmod_reg) begin
                        if (reg_wait)   CS_usr <= CS ;
			else if (CS_enable) CS_usr <= mdw_pre[3:0] ;
                end
        end

        //synopsys async_set_reset "resb"
        always @(posedge baseck or negedge resb) begin
                if (!resb)              CS_sv <= 4'h0 ;
                else if (cpuen && sel_svmod_reg) begin
                        if (reg_wait)   CS_sv <= CS ;
			else if (CS_enable) CS_sv <= mdw_pre[3:0] ;
                end
        end
//

/*------------------------------------------------------------------------------*/
/* �ץ��å��⡼�ɥ���ȥ���쥸���� �Уͣ�					*/
/*------------------------------------------------------------------------------*/
/*   �ң��Ͷ��֤إߥ顼����ե�å��������֤����򤹤롣			*/
/*------------------------------------------------------------------------------*/

// MAA�����ʤ�00000H��0FFFFH��F0000H��FFFFFH�إߥ顼���롣
// MAA�����ʤ�10000H��1FFFFH��F0000H��FFFFFH�إߥ顼���롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)
			MAA <= 1'b0;
		else if (cpuen) begin
			if (reg_wait)	MAA <= MAA ;
			else if (pselcpu && cpuwr) begin
				casex (vpa)
					4'he : MAA <= mdw_pre[0] ;
					default	: MAA <= MAA ;
				endcase
			end
		end
	end

/*------------------------------------------------------------------------------*/
/* �꡼�ɡ��饤�ȥ��͡��֥뿮��							*/
/*------------------------------------------------------------------------------*/
/*   �ǡ�������ڤӣӣƣҶ��֤ؤΥ꡼�ɡ��饤�ȥ��͡��֥뿮����������롣	*/
/*------------------------------------------------------------------------------*/

// �ǡ������������򼨤����档RAM�ؤΥե��å����������ȶ��̤���٤˻��Ѥ��롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)		mem_access <= 1'b0 ;
		else if (cpuen) begin
					mem_access <= dec_cpuwr_enable | dec_cpurd_enable ;
		end
	end

// �ǥ���������Υ꡼�ɡ��饤�ȿ���������쥸������
// �ϥ�����ȯ������BTCLR�������Ω������ť����������ɤ�����cpuwr_pre��cpurd_pre�ϣ��ˤʤ롣
// RAM�ե��å����̿�����ɤ߾��֤ΤȤ���cpuwr_pre�ϣ��Ȥʤꡢ�դ�̿�����ɤ߾��֤�cpurd_pre�ϣ��Ȥʤ롣
// �ޤ�RAM�ե��å����cpurd_pre�ϥ饤�ȥ����������ˤϣ��Ȥʤ롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) begin
			cpuwr_pre <= 1'b0 ;
			cpurd_pre <= 1'b0 ;
		end
		else if (cpuen) begin
// ʬ���������Ω���ˡ��꡼�ɡ��饤�ȥ��ȥ��֤�Ω��������Τϡ�
// ���ꥢ��������Ȥ�ʤ�ʬ��̿��Τߡ�
			if (data_hazard_flg || (stage_cut && dec_ma_enable)) begin
				cpuwr_pre <= 1'b0 ;
				cpurd_pre <= 1'b0 ;
			end
			else if (fchiram) begin
				cpuwr_pre <= dec_cpuwr_enable & ~pa_st2 ;
				cpurd_pre <= dec_cpurd_enable | ~dec_cpuwr_enable | pa_st2 ;
			end
			else begin
				cpuwr_pre <= dec_cpuwr_enable ;
				cpurd_pre <= dec_cpurd_enable ;
			end
		end
	end

// ����ؤΥ饤�ȡ��꡼�ɥ��ȥ��ֿ��档
// DMAž�����dmawr��dmard�����줾�����򤵤�롣
	assign cpuwr_reg = ~sp_sfr_en & cpuwr_pre;
	assign cpuwr = (waitdma) ? dmawr : ~sp_sfr_en & cpuwr_pre ;
	assign cpurd = (waitdma) ? dmard : cpurd_pre ;

// RAM�ե��å���˥���ؤΥ꡼�ɥ���������ȯ��������磱�Ȥʤ롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)			fchiram_cpurd <= 1'b0 ;
		else if (cpuen) begin
			if (fchiram)		fchiram_cpurd <= dec_cpurd_enable ;
			else			fchiram_cpurd <= 1'b0 ;
		end
	end

/*------------------------------------------------------------------------------*/
/* ���Ƚ�꿮��									*/
/*------------------------------------------------------------------------------*/
/*   ���ʬ��̿��¹Ի��˾��Ƚ���Ԥʤ���					*/
/*------------------------------------------------------------------------------*/

// C�ޤ���Z�ˤ��ʬ�����Ƚ�꿮�档
// �����������Ȥ�HIGH���򣱥���å�������Ф���
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) 		stage_cut_ifbr <= 1'b0 ;
		else if (cpuen) begin
			if (pc_wait_flg)	stage_cut_ifbr <= stage_cut_ifbr ;
			else			stage_cut_ifbr <= dec_stage_cut_ifbr ;
		end
	end

// ʬ�����Ƚ�꿮�档�����������Ȥ�HIGH���򣱥���å�������Ф���
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) 		stage_cut_brtf <= 1'b0 ;
		else if (cpuen) begin
			if (pc_wait_flg)	stage_cut_brtf <= stage_cut_brtf ;
			else			stage_cut_brtf <= dec_stage_cut_brtf ;
		end
	end

// ʬ��̿��ˤ��PSW���������ǤΥ������Ȥ򤳤ο�����ޤ��롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) 		wait_block_brtf <= 1'b0 ;
		else if (cpuen) begin
			if (pc_wait_flg)	wait_block_brtf <= wait_block_brtf ;
			else			wait_block_brtf <= stage_cut_brtf ;
		end
	end

// ���ʬ��̿��¹Ի��ˣ��Ȥʤ롣
	assign stage_cut_br = stage_cut_ifbr | stage_cut_brtf ;

// RAM�ե��å���ξ��Ƚ��ϣ�����å��٤��Τǡ�Ƚ���̤��ݻ����Ƥ�����
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) 		stage_cut_alu <= 1'b0 ;
		else if (cpuen) begin
			if (pc_wait_flg)	stage_cut_alu <= stage_cut_alu ;
			else if (fchiram)	stage_cut_alu <= ~buf0[0] ;
			else			stage_cut_alu <= ~aluout[0] ;
		end
	end

// Ƚ���郎ZȽ��ξ��ifbr_zero����CȽ��ξ�磰�Ȥʤ롣
// �ޤ���Ƚ���郎��Ƚ��ξ��ifbr_not��������Ƚ��ξ�磰�Ȥʤ롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) begin
				ifbr_not <= 1'b0 ;
				ifbr_zero <= 1'b0 ;
				ifbr_ht <= 1'b0 ;
		end
		else if (cpuen) begin
			if (pc_wait_flg) begin
				ifbr_not <= ifbr_not ;
				ifbr_zero <= ifbr_zero ;
				ifbr_ht <= ifbr_ht ;
			end
			else begin
				ifbr_not <= dec_ifbr_not ;
				ifbr_zero <= dec_ifbr_zero ;
				ifbr_ht <= dec_ifbr_ht ;
			end
		end
	end

// ʬ����郎����Ω�ξ�磱�Ȥʤꡢʬ��̿��μ¹Ԥ���Ū�˽�λ���롣
// BRT/F/TCLR���ϥ��ԡ��ɤ�����ǡ�Ƚ��ӥåȤ��ݻ��Хåե��˳�Ǽ���Ƥ�����
	always @(fchiram or stage_cut_ifbr or stage_cut_brtf or ifbr_not or ifbr_zero or ifbr_ht or
		 stage_cut_alu or CY or Z or buf0) begin
		if (stage_cut_ifbr) begin
			casex ({ifbr_not,ifbr_zero,ifbr_ht})
				3'b000	: stage_cut = ~CY ;
				3'b100	: stage_cut = CY ;
				3'b010	: stage_cut = ~Z ;
				3'b110	: stage_cut = Z ;
				3'b001	: stage_cut = (Z | CY) ;
				3'b101	: stage_cut = ~(Z | CY) ;
				default	: stage_cut = 1'b0 ;
			endcase
		end
		else if (stage_cut_brtf) begin
			if (fchiram)		stage_cut = stage_cut_alu ;
			else			stage_cut = ~buf0[0] ;
		end
		else				stage_cut = 1'b0 ;
	end

/*------------------------------------------------------------------------------*/
/* �����åץե饰								*/
/*------------------------------------------------------------------------------*/
/*   �����åץե饰���������롣							*/
/*------------------------------------------------------------------------------*/

// SKIP̿��¹Ի��˳������׵����α���뤿��ο��档
	assign skp_block = dec_skc | dec_sknc | dec_skz | dec_sknz | dec_skh | dec_sknh ;

// �����å�Ƚ�꿮�档�����å�̿���Ƚ��������椹�롣
// ������������ȯ�����ޤ������ɤ߾��֤Ǥ��ݻ�����롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) begin
			skip_c  <= 1'b0 ;
			skip_nc <= 1'b0 ;
			skip_z  <= 1'b0 ;
			skip_nz <= 1'b0 ;
			skip_h  <= 1'b0 ;
			skip_nh <= 1'b0 ;
		end
		else if (cpuen) begin
			if (pc_wait_flg || pa_st2) begin
				skip_c  <= skip_c ;
				skip_nc <= skip_nc ;
				skip_z  <= skip_z ;
				skip_nz <= skip_nz ;
				skip_h  <= skip_h ;
				skip_nh <= skip_nh ;
			end
			else begin
				skip_c  <= dec_skc ;
				skip_nc <= dec_sknc ;
				skip_z  <= dec_skz ;
				skip_nz <= dec_sknz ;
				skip_h  <= dec_skh ;
				skip_nh <= dec_sknh ;
			end
		end
	end

// �����å��о�̿�᤬PREFIX̿����ä�����skpack��̿��ʬȯ�Ԥ��롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) 			prefix_skp <= 1'b0 ;
		else if (cpuen) begin
			if (pc_wait_flg)	prefix_skp <= prefix_skp ;
			else if (skpack && !(fchiram_skp || romrd_skp) && (ID_stage0 == 8'h11))
						prefix_skp <= 1'b1 ;
			else			prefix_skp <= 1'b0 ;
		end
	end

// �����å׼¹ԥե饰�������å׾������򤷡��ǥ�������skpack���Ϥ���
// FLASH�ե��å����FLASH�ؤΥǡ�������������ȯ���������ȡ�
// RAM�ե��å����RAM����������ȯ��������硢���פ�̿��μ¹Ԥ��ɤ����ᤳ�ο�����Ѥ��롣
	always @(skip_c or skip_nc or skip_z or skip_nz or skip_h or skip_nh or
		 CY or Z or prefix_skp or fchiram_skp or romrd_skp) begin
		if (skip_c)				skpack = CY ;
		else if (skip_nc)			skpack = ~CY ;
		else if (skip_z)			skpack = Z ;
		else if (skip_nz)			skpack = ~Z ;
		else if (skip_h)			skpack = ~(CY | Z) ;
		else if (skip_nh)			skpack = (CY | Z) ;
		else if (prefix_skp)			skpack = 1'b1 ;
		else if (fchiram_skp || romrd_skp)	skpack = 1'b1 ;
		else					skpack = 1'b0 ;
	end

// �����å׾�郎��Ω�����о�̿�᤬�����åפ��줿����ɽ�����档
	assign skipexe = skpack & ~fchiram_skp & ~romrd_skp ;

/*------------------------------------------------------------------------------*/
/* �£ã�����									*/
/*------------------------------------------------------------------------------*/
/*   �£ã������ǡ���������꡼�����ǡ������������롣				*/
/*------------------------------------------------------------------------------*/

// �黻��̤β��̣��ӥåȤ�������ɬ�פʾ�磱�Ȥʤ롣
	assign	bcdadj_low = A[3] & (A[2] | A[1]) ;

// �黻��̤���������ɬ�פʾ��ϡ����Ȥʤ롣
	assign	bcdadj_flg[0] = AC | bcdadj_low ;
	assign	bcdadj_flg[1] = CY | (A[7] & (A[6] | A[5] | (A[4] & bcdadj_low))) ;

// BCDADJ�쥸�������ɤߤ����ͤϡ�A�쥸���������������͡�
	assign	BCDADJ = bcdadj_flg ;

endmodule


/*------------------------------------------------------------------------------*/
/* ���������黻��˥å�								*/
/*------------------------------------------------------------------------------*/
/*   ���������黻��¹Ԥ��롣							*/
/*------------------------------------------------------------------------------*/
/* Ver2.0  �ӥå�̿�ᡢ���ե�̿������ƺ����					*/
/*------------------------------------------------------------------------------*/
module QLK0RCPUEVA0V3_EXE(
		aluin10, aluin11, aluin20, aluin21, CY,
		dec_alu_add, dec_alu_sub, dec_alu_and, dec_alu_or, dec_alu_exor,
		dec_alu_carry, dec_word_access,
		exeout, acout, cyout
		);

	input	[7:0]	aluin10, aluin11, aluin20, aluin21;
	input		dec_alu_add, dec_alu_sub, dec_alu_and, dec_alu_or, dec_alu_exor;
	input		dec_alu_carry, dec_word_access;
	input		CY;

	output	[15:0]	exeout;
	output		acout, cyout;

	reg	[15:0]	exeout;
	reg		acout, cyout;
	reg		cy_byte, cy_word;

// ALU�ε�ǽ�����򤷡��黻��¹Ԥ��롣
// �������̾��Τ��ᡢ���Ƥ�̿�᤬������ʬ���̲᤹�롣
	always @(aluin10 or aluin11 or aluin20 or aluin21 or CY or
		 dec_alu_add or dec_alu_sub or dec_alu_and or dec_alu_or or dec_alu_exor or
		 dec_alu_carry or dec_word_access) begin
		if (dec_alu_add) begin //ADD
			{acout,   exeout[3:0]}  = {1'b0,aluin10[3:0]} + {1'b0,aluin20[3:0]} + (CY & dec_alu_carry) ;
			{cy_byte, exeout[7:4]}  = {1'b0,aluin10[7:4]} + {1'b0,aluin20[7:4]} + acout ;
			{cy_word, exeout[15:8]} = {1'b0,aluin11} + {1'b0,aluin21} + cy_byte ;
			if (dec_word_access) cyout = cy_word ;
			else cyout = cy_byte ;
		end
		else if (dec_alu_sub) begin //SUB
			{acout,   exeout[3:0]}  = {1'b0,aluin10[3:0]} - {1'b0,aluin20[3:0]} - (CY & dec_alu_carry) ;
			{cy_byte, exeout[7:4]}  = {1'b0,aluin10[7:4]} - {1'b0,aluin20[7:4]} - acout ;
			{cy_word, exeout[15:8]} = {1'b0,aluin11} - {1'b0,aluin21} - cy_byte ;
			if (dec_word_access) cyout = cy_word ;
			else cyout = cy_byte ;
		end
		else if (dec_alu_and) begin //AND
			exeout[15:8] = 8'h00 ;
			exeout[7:0] = aluin10 & aluin20 ;
			acout = 1'b0 ;
			cyout = 1'b0 ;
		end
		else if (dec_alu_or) begin //OR
			exeout[15:8] = 8'h00 ;
			exeout[7:0] = aluin10 | aluin20 ;
			acout = 1'b0 ;
			cyout = 1'b0 ;
		end
		else if (dec_alu_exor) begin //EXOR
			exeout[15:8] = 8'h00 ;
			exeout[7:0] = aluin10 ^ aluin20 ;
			acout = 1'b0 ;
			cyout = 1'b0 ;
		end
		else begin  //MOV
			exeout = {aluin21,aluin20} ;
			acout = 1'b0 ;
			cyout = 1'b0 ;
		end
	end

endmodule

/*------------------------------------------------------------------------------*/
/* ���������黻��˥å�                                                         */
/*------------------------------------------------------------------------------*/
/* Ver2.0  ���������黻��¹Ԥ��롣						*/
/*------------------------------------------------------------------------------*/
module QLK0RCPUEVA0V3_EXE2(
                bitshin10, bitshin20, bitshin21, CY,
                dec_alu_andbit, dec_alu_orbit, dec_alu_exorbit,
                dec_alu_ror, dec_alu_rol, dec_alu_shr, dec_alu_shl, dec_alu_sar,
                dec_alu_carry, MEM_stage0h, dec_word_access,
                bitshout, cyout
                );

        input   [7:0]   bitshin10, bitshin20, bitshin21;
        input   [3:0]   MEM_stage0h;
        input           dec_alu_andbit, dec_alu_orbit, dec_alu_exorbit;
        input           dec_alu_ror, dec_alu_rol, dec_alu_shr, dec_alu_shl, dec_alu_sar;
        input           dec_alu_carry, dec_word_access;
        input           CY;

        output  [15:0]  bitshout;
        output          cyout;

        reg     [15:0]  bitshout;
        reg             cyout;
        reg             cy_byte, cy_word;

// ALU�ε�ǽ�����򤷡��黻��¹Ԥ��롣
// �������̾��Τ��ᡢ���Ƥ�̿�᤬������ʬ���̲᤹�롣
// ���ե�̿��ϥ��ڥ�������˥��ե����������ޤ�Ƥ���Τǡ�MEM���ơ����쥸�����Υǡ������ɤ߹��ࡣ
        always @(bitshin10 or bitshin20 or bitshin21 or CY or
                 dec_alu_andbit or dec_alu_orbit or dec_alu_exorbit or
                 dec_alu_ror or dec_alu_rol or dec_alu_shr or dec_alu_shl or dec_alu_sar or
                 dec_alu_carry or MEM_stage0h or dec_word_access) begin
                if (dec_alu_andbit) begin //AND1,CLR1
                        bitshout[15:8] = 8'h00 ;
                        bitshout[7:0] = bitshin10 & bitshin20 ;
                        cyout = 1'b0 ;
                end
                else if (dec_alu_orbit) begin //OR1,SET1
                        bitshout[15:8] = 8'h00 ;
                        bitshout[7:0] = bitshin10 | bitshin20 ;
                        cyout = 1'b0 ;
                end
                else if (dec_alu_exorbit) begin //EXOR1,NOT1
                        bitshout[15:8] = 8'h00 ;
                        bitshout[7:0] = bitshin10 ^ bitshin20 ;
                        cyout = 1'b0 ;
                end
                else if (dec_alu_ror) begin //ROR
                        bitshout[15:8] = 8'h00 ;
                        bitshout[7]   = (dec_alu_carry) ? CY : bitshin20[0] ;
                        bitshout[6:0] = bitshin20[7:1] ;
                        cyout = bitshin20[0] ;
                end
                else if (dec_alu_rol) begin //ROL
                        if (dec_word_access) begin
                                bitshout[15:1] = {bitshin21[6:0],bitshin20[7:0]} ;
                                bitshout[0] = (dec_alu_carry) ? CY : bitshin21[7] ;
                                cyout = bitshin21[7] ;
                        end
                        else begin
                                bitshout[15:8] = 8'h00 ;
                                bitshout[0]   = (dec_alu_carry) ? CY : bitshin20[7] ;
                                bitshout[7:1] = bitshin20[6:0] ;
                                cyout = bitshin20[7] ;
                        end
                end
                else if (dec_alu_shr) begin //SHR
                        casex ({MEM_stage0h,dec_word_access})
                                ({4'h1,1'b0}) : {bitshout,cyout} = {8'h00,1'b0,bitshin20[7:1],bitshin20[0]} ;
                                ({4'h2,1'b0}) : {bitshout,cyout} = {8'h00,2'b0,bitshin20[7:2],bitshin20[1]} ;
                                ({4'h3,1'b0}) : {bitshout,cyout} = {8'h00,3'b0,bitshin20[7:3],bitshin20[2]} ;
                                ({4'h4,1'b0}) : {bitshout,cyout} = {8'h00,4'b0,bitshin20[7:4],bitshin20[3]} ;
                                ({4'h5,1'b0}) : {bitshout,cyout} = {8'h00,5'b0,bitshin20[7:5],bitshin20[4]} ;
                                ({4'h6,1'b0}) : {bitshout,cyout} = {8'h00,6'b0,bitshin20[7:6],bitshin20[5]} ;
                                ({4'h7,1'b0}) : {bitshout,cyout} = {8'h00,7'b0,bitshin20[7],bitshin20[6]} ;
                                ({4'h0,1'b1}) : {bitshout,cyout} = { bitshin21[7:0],bitshin20[7:0],1'b0} ;
                                ({4'h1,1'b1}) : {bitshout,cyout} = { 1'b0,bitshin21[7:0],bitshin20[7:1],bitshin20[0]} ;
                                ({4'h2,1'b1}) : {bitshout,cyout} = { 2'b0,bitshin21[7:0],bitshin20[7:2],bitshin20[1]} ;
                                ({4'h3,1'b1}) : {bitshout,cyout} = { 3'b0,bitshin21[7:0],bitshin20[7:3],bitshin20[2]} ;
                                ({4'h4,1'b1}) : {bitshout,cyout} = { 4'b0,bitshin21[7:0],bitshin20[7:4],bitshin20[3]} ;
                                ({4'h5,1'b1}) : {bitshout,cyout} = { 5'b0,bitshin21[7:0],bitshin20[7:5],bitshin20[4]} ;
                                ({4'h6,1'b1}) : {bitshout,cyout} = { 6'b0,bitshin21[7:0],bitshin20[7:6],bitshin20[5]} ;
                                ({4'h7,1'b1}) : {bitshout,cyout} = { 7'b0,bitshin21[7:0],bitshin20[7],bitshin20[6]} ;
                                ({4'h8,1'b1}) : {bitshout,cyout} = { 8'b0,bitshin21[7:0],bitshin20[7]} ;
                                ({4'h9,1'b1}) : {bitshout,cyout} = { 9'b0,bitshin21[7:1],bitshin21[0]} ;
                                ({4'ha,1'b1}) : {bitshout,cyout} = {10'b0,bitshin21[7:2],bitshin21[1]} ;
                                ({4'hb,1'b1}) : {bitshout,cyout} = {11'b0,bitshin21[7:3],bitshin21[2]} ;
                                ({4'hc,1'b1}) : {bitshout,cyout} = {12'b0,bitshin21[7:4],bitshin21[3]} ;
                                ({4'hd,1'b1}) : {bitshout,cyout} = {13'b0,bitshin21[7:5],bitshin21[4]} ;
                                ({4'he,1'b1}) : {bitshout,cyout} = {14'b0,bitshin21[7:6],bitshin21[5]} ;
                                ({4'hf,1'b1}) : {bitshout,cyout} = {15'b0,bitshin21[7],bitshin21[6]} ;
                                default : {bitshout,cyout} = {8'h00,bitshin20,1'b0} ;
                        endcase
                end
                else if (dec_alu_shl) begin //SHL
                        casex ({MEM_stage0h,dec_word_access})
                                ({4'h1,1'b0}) : {bitshout,cyout} = {8'h00,bitshin20[6:0],1'b0,bitshin20[7]} ;
                                ({4'h2,1'b0}) : {bitshout,cyout} = {8'h00,bitshin20[5:0],2'b0,bitshin20[6]} ;
                                ({4'h3,1'b0}) : {bitshout,cyout} = {8'h00,bitshin20[4:0],3'b0,bitshin20[5]} ;
                                ({4'h4,1'b0}) : {bitshout,cyout} = {8'h00,bitshin20[3:0],4'b0,bitshin20[4]} ;
                                ({4'h5,1'b0}) : {bitshout,cyout} = {8'h00,bitshin20[2:0],5'b0,bitshin20[3]} ;
                                ({4'h6,1'b0}) : {bitshout,cyout} = {8'h00,bitshin20[1:0],6'b0,bitshin20[2]} ;
                                ({4'h7,1'b0}) : {bitshout,cyout} = {8'h00,bitshin20[0],7'b0,bitshin20[1]} ;
                                ({4'h0,1'b1}) : {bitshout,cyout} = {bitshin21[7:0],bitshin20[7:0],1'b0} ;
                                ({4'h1,1'b1}) : {bitshout,cyout} = {bitshin21[6:0],bitshin20[7:0],1'b0,bitshin21[7]} ;
                                ({4'h2,1'b1}) : {bitshout,cyout} = {bitshin21[5:0],bitshin20[7:0],2'b0,bitshin21[6]} ;
                                ({4'h3,1'b1}) : {bitshout,cyout} = {bitshin21[4:0],bitshin20[7:0],3'b0,bitshin21[5]} ;
                                ({4'h4,1'b1}) : {bitshout,cyout} = {bitshin21[3:0],bitshin20[7:0],4'b0,bitshin21[4]} ;
                                ({4'h5,1'b1}) : {bitshout,cyout} = {bitshin21[2:0],bitshin20[7:0],5'b0,bitshin21[3]} ;
                                ({4'h6,1'b1}) : {bitshout,cyout} = {bitshin21[1:0],bitshin20[7:0],6'b0,bitshin21[2]} ;
                                ({4'h7,1'b1}) : {bitshout,cyout} = {bitshin21[0],bitshin20[7:0],7'b0,bitshin21[1]} ;
                                ({4'h8,1'b1}) : {bitshout,cyout} = {bitshin20[7:0], 8'b0,bitshin21[0]} ;
                                ({4'h9,1'b1}) : {bitshout,cyout} = {bitshin20[6:0], 9'b0,bitshin20[7]} ;
                                ({4'ha,1'b1}) : {bitshout,cyout} = {bitshin20[5:0],10'b0,bitshin20[6]} ;
                                ({4'hb,1'b1}) : {bitshout,cyout} = {bitshin20[4:0],11'b0,bitshin20[5]} ;
                                ({4'hc,1'b1}) : {bitshout,cyout} = {bitshin20[3:0],12'b0,bitshin20[4]} ;
                                ({4'hd,1'b1}) : {bitshout,cyout} = {bitshin20[2:0],13'b0,bitshin20[3]} ;
                                ({4'he,1'b1}) : {bitshout,cyout} = {bitshin20[1:0],14'b0,bitshin20[2]} ;
                                ({4'hf,1'b1}) : {bitshout,cyout} = {bitshin20[0],15'b0,bitshin20[1]} ;
                                default : {bitshout,cyout} = {8'h00,bitshin20,1'b0} ;
                        endcase
                end
                else if (dec_alu_sar) begin //SAR
                        casex ({MEM_stage0h,dec_word_access})
                                ({4'h1,1'b0}) : {bitshout,cyout} = {8'h00,bitshin20[7],bitshin20[7:1],bitshin20[0]} ;
                                ({4'h2,1'b0}) : {bitshout,cyout} = {8'h00,{2{bitshin20[7]}},bitshin20[7:2],bitshin20[1]} ;
                                ({4'h3,1'b0}) : {bitshout,cyout} = {8'h00,{3{bitshin20[7]}},bitshin20[7:3],bitshin20[2]} ;
                                ({4'h4,1'b0}) : {bitshout,cyout} = {8'h00,{4{bitshin20[7]}},bitshin20[7:4],bitshin20[3]} ;
                                ({4'h5,1'b0}) : {bitshout,cyout} = {8'h00,{5{bitshin20[7]}},bitshin20[7:5],bitshin20[4]} ;
                                ({4'h6,1'b0}) : {bitshout,cyout} = {8'h00,{6{bitshin20[7]}},bitshin20[7:6],bitshin20[5]} ;
                                ({4'h7,1'b0}) : {bitshout,cyout} = {8'h00,{7{bitshin20[7]}},bitshin20[7],bitshin20[6]} ;
                                ({4'h0,1'b1}) : {bitshout,cyout} = {bitshin21[7:0],bitshin20[7:0],1'b0} ;
                                ({4'h1,1'b1}) : {bitshout,cyout} = {bitshin21[7],bitshin21[7:0],bitshin20[7:1],bitshin20[0]} ;
                                ({4'h2,1'b1}) : {bitshout,cyout} = {{ 2{bitshin21[7]}},bitshin21[7:0],bitshin20[7:2],bitshin20[1]} ;
                                ({4'h3,1'b1}) : {bitshout,cyout} = {{ 3{bitshin21[7]}},bitshin21[7:0],bitshin20[7:3],bitshin20[2]} ;
                                ({4'h4,1'b1}) : {bitshout,cyout} = {{ 4{bitshin21[7]}},bitshin21[7:0],bitshin20[7:4],bitshin20[3]} ;
                                ({4'h5,1'b1}) : {bitshout,cyout} = {{ 5{bitshin21[7]}},bitshin21[7:0],bitshin20[7:5],bitshin20[4]} ;
                                ({4'h6,1'b1}) : {bitshout,cyout} = {{ 6{bitshin21[7]}},bitshin21[7:0],bitshin20[7:6],bitshin20[5]} ;
                                ({4'h7,1'b1}) : {bitshout,cyout} = {{ 7{bitshin21[7]}},bitshin21[7:0],bitshin20[7],bitshin20[6]} ;
                                ({4'h8,1'b1}) : {bitshout,cyout} = {{ 8{bitshin21[7]}},bitshin21[7:0],bitshin20[7]} ;
                                ({4'h9,1'b1}) : {bitshout,cyout} = {{ 9{bitshin21[7]}},bitshin21[7:1],bitshin21[0]} ;
                                ({4'ha,1'b1}) : {bitshout,cyout} = {{10{bitshin21[7]}},bitshin21[7:2],bitshin21[1]} ;
                                ({4'hb,1'b1}) : {bitshout,cyout} = {{11{bitshin21[7]}},bitshin21[7:3],bitshin21[2]} ;
                                ({4'hc,1'b1}) : {bitshout,cyout} = {{12{bitshin21[7]}},bitshin21[7:4],bitshin21[3]} ;
                                ({4'hd,1'b1}) : {bitshout,cyout} = {{13{bitshin21[7]}},bitshin21[7:5],bitshin21[4]} ;
                                ({4'he,1'b1}) : {bitshout,cyout} = {{14{bitshin21[7]}},bitshin21[7:6],bitshin21[5]} ;
                                ({4'hf,1'b1}) : {bitshout,cyout} = {{15{bitshin21[7]}},bitshin21[7],bitshin21[6]} ;
                                default : {bitshout,cyout} = {8'h00,bitshin20,1'b0} ;
                        endcase
                end
//              else if (dec_alu_mulu) begin //MULU teg3
//                      bitshout = bitshin10 * bitshin20 ;
//                      acout = 1'b0 ;
//                      cyout = 1'b0 ;
//              end
                else begin  //MOV
                        bitshout = {bitshin21,bitshin20} ;
                        cyout = 1'b0 ;
                end
        end

endmodule

/********************************************************************************/
/* K0R EVA CLK Block                                                           	*/
/*                                                          Made K.Tanaka       */
/********************************************************************************/
/* Ver1.00  New                                                                 */
/* Ver1.50  Add stbst                                 2007.07.02 K.Tanaka       */
/********************************************************************************/
module QLK0RCPUEVA0V3_CLK(
	mdr, imdr, pselcpu, pselbcd, slreg, rga, vpa,
	dec_set_buf_retadr, dec_set_buf_intr,
	dec_halt, dec_stop, stben, pc_wait_flg, stby_wait_flg, cpurd, wdop,
	intdbg, intnmi, intrq3, intrq2, intrq1, intrq0,
	SP, PSW, CS, ES, MAA, BCDADJ,
	A_bank0, X_bank0, B_bank0, C_bank0, D_bank0, E_bank0, H_bank0, L_bank0,
	A_bank1, X_bank1, B_bank1, C_bank1, D_bank1, E_bank1, H_bank1, L_bank1,
	A_bank2, X_bank2, B_bank2, C_bank2, D_bank2, E_bank2, H_bank2, L_bank2,
	A_bank3, X_bank3, B_bank3, C_bank3, D_bank3, E_bank3, H_bank3, L_bank3,
	INT_wait, wait2ndsfr, sl2ndwait_pre, waitdma, waitint, dmarq, dopen, dmaack,
	waitfl, waitmod, waitexm, dmaen, dmawait, ocdwait, pswlock,
	exmmsk, flmask, hltst, stpst, stbst,
// for EVA
        SP_usr, SP_sv, svmod, alt1,
        svi,
        waitfl2, icewaitmem,
        cpumask,
//
	cpustart, cpuen, pswen, baseck, resb, scanmode,
	sldfwait_pre, waitdflash,
	RVEON, crchlten
	);

	output	[15:0]	imdr;
	output		cpuen, pswen;
	output		pswlock;
	output		waitint, waitdma;
	output		dmawait, dmaack;
	output		ocdwait;
	output		stben;
	output		exmmsk;
	output		flmask;
	output		hltst, stpst;
	output		stbst;		// add v1.50 2007.07.02 K.Tanaka

// for EVA
        output          cpumask;
//

	input	[15:0]	mdr;
	input		pselcpu, pselbcd;
	input		slreg;
	input		rga;
	input	[3:0]	vpa;
	input		dec_set_buf_retadr, dec_set_buf_intr;
	input		dec_halt, dec_stop;
	input		pc_wait_flg, stby_wait_flg;
	input		cpurd, wdop;
	input	[14:0]	SP;
	input	[7:0]	PSW;
	input	[3:0]	CS, ES;
	input		MAA;
	input	[1:0]	BCDADJ;
	input	[7:0]	A_bank0,X_bank0,B_bank0,C_bank0,D_bank0,E_bank0,H_bank0,L_bank0;
	input	[7:0]	A_bank1,X_bank1,B_bank1,C_bank1,D_bank1,E_bank1,H_bank1,L_bank1;
	input	[7:0]	A_bank2,X_bank2,B_bank2,C_bank2,D_bank2,E_bank2,H_bank2,L_bank2;
	input	[7:0]	A_bank3,X_bank3,B_bank3,C_bank3,D_bank3,E_bank3,H_bank3,L_bank3;
	input		intdbg, intnmi, intrq3, intrq2, intrq1, intrq0;
	input		INT_wait, wait2ndsfr, sl2ndwait_pre;
	input		waitfl, waitmod, waitexm;
	input		dmarq, dopen;
	input		dmaen;
	input		cpustart;
	input		baseck, resb;
	input		scanmode;
	input		sldfwait_pre;
	input		waitdflash;
	input		RVEON;
	input		crchlten;
// for EVA
        input   [14:0]  SP_usr, SP_sv;
        input           svmod;
        input           alt1;
        input           svi;
        input           waitfl2, icewaitmem;
//

	wire		stby, stben;
	wire		cpuen_pre;
	wire		flmask_pre;
	wire		waitdma;

// for EVA
        wire    [14:0]  SP_rd;
//

	reg	[15:0]	cpumdr;
	reg	[1:0]	wait_cnt;
	reg		waitint;
	reg		dmaack_pre;
	reg		DMA_read, DMA_write;

/*------------------------------------------------------------------------------*/
/* �ãУե��͡��֥�								*/
/*------------------------------------------------------------------------------*/
/*   �ȣ��̣ԡ��ӣԣϣ�̿��¹Ի��ȳ�����������ȯ�����˥���å�����ߤ����롣	*/
/*------------------------------------------------------------------------------*/

// CPU�����������Ȥǡ�CPU��ǥ����������򥫥���Ȥ�����Υ����󥿡�
// INT̿���INT�ޥ����SFR��PSW�ؤν񤭹��߶������򤹤륦�����Ȥǥ�����ȥ��åס�
// DMAž���桢�ޤ��ϳ�������������ϥ�����ȥ��åפ��ƤϤ����ʤ���
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb) begin
			wait_cnt <= 2'h0 ;
		end
		else if (waitdma || waitexm || wait2ndsfr || waitdflash || waitfl || waitmod) begin
			wait_cnt <= wait_cnt ;
		end
		else if (waitint) begin
			wait_cnt <= wait_cnt + 2'h1 ;
		end
		else begin
			wait_cnt <= 2'h0 ;
		end
	end

// ����������WAITINT��������å��������ȤʤΤǡ�
// �������ȥ�����ȣ���Ω�������롣
	always @(INT_wait or wait_cnt) begin
		if (INT_wait)
			if (wait_cnt == 2'h2)	waitint = 1'b0 ;
			else			waitint = 1'b1 ;
		else				waitint = 1'b0 ;
	end

// dmarq������դ�������Ω���夬�롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)			dmaack_pre <= 1'b0 ;
		else if (dmaen) begin
			if (dmawait)		dmaack_pre <= dmaack_pre ;
			else if (dmaack_pre)	dmaack_pre <= 1'b0 ;
			else			dmaack_pre <= dopen & dmarq ;
		end
	end

// CALL�ʤ�ID���ơ������ݻ��Хåե�����Ѥ���̿�ᡢ̿��ˤ��WAIT
// �Υ�ޥ����֥�������׵�ȯ����DMAACK��ޥ������롣
// for EVA
//	assign dmaack = dmaack_pre & ~(dec_set_buf_retadr | dec_set_buf_intr) & ~waitint & ~sl2ndwait_pre & ~(intdbg | intnmi) ;
	assign dmaack = dmaack_pre & ~(dec_set_buf_retadr | dec_set_buf_intr) & ~waitint & ~sl2ndwait_pre & ~sldfwait_pre & ~(intdbg | intnmi | svi) ;
//

// DMA�Υ꡼�ɥ��������ɽ�����档
// DMA�����դ����ˣ��Ȥʤ롣
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)		DMA_read <= 1'b0 ;
		else if (dmaen) begin
			if (dmawait)	DMA_read <= DMA_read ;
			else		DMA_read <= dmaack ;
		end
	end

// DMA�Υ饤�ȥ��������ɽ�����档
// DMAž����Υ������ȿ���򣱥���å���Ф���
	//synopsys async_set_reset "resb"
	always @(posedge baseck or negedge resb) begin
		if (!resb)		DMA_write <= 1'b0 ;
		else if (dmaen) begin
			if (dmawait)	DMA_write <= DMA_write ;
			else		DMA_write <= DMA_read ;
		end
	end

// DMAž����Υ������ȿ��档
	assign waitdma = DMA_read | DMA_write ;

// DMAž�����slexm�����ޥ������Х����������ȯ�Ԥ��Ԥ�����٤ο��档
// ����������쥸�����Υ饤�ȥ��������ˤ�륦�����ȤǤ�slexm��ޥ������롣
	assign exmmsk = DMA_read | (DMA_write & dmawait) | waitint ;

// WAITINTȯ������PSW������ư�������档
	assign pswen = waitint & (wait_cnt == 2'b00) & ~waitdma ;

// PSW���������Υ������Ȥˤ����ơ�PSW�ι����Ϻǽ�Σ�����å��Τߡ�
// ����ʳ��δ��֤Ϥ��ο�����ݻ����롣
	assign pswlock = wait_cnt[1] | wait_cnt[0] ;

// �������׵᤬�����磱�Ȥʤ롣���λ���������Х����֤ˤ�����ʤ���
// for EVA
//	assign stben = intdbg | intnmi | intrq3 | intrq2 | intrq1 | intrq0 ;
        assign stben = intdbg | intnmi | intrq3 | intrq2 | intrq1 | intrq0 | crchlten | svi ;
//

// HALT/STOP̿�᤬�¹Ԥ��줿�Ȥ����Ȥʤ롣
	assign stbst = dec_halt | dec_stop ;

// HALT̿��STOP̿��¹Ի��ˣ��Ȥʤ롣�������׵᤬������ϣ���
// RAM�ե��å����̿��ե��å�����(pc_wait_flg)��HALT/STOP������ʤ���
/*------------------------------------------------------------------------------*/
/* Ver2.0  SLFLASH�Υ��ԡ��ɥ��åפΰ١�pc_wait_flg���ѹ����롣			*/
/*��������������RAM�ե��å���HALT�ǻߤޤä��ݤˡ��ߤޤ��꤬RAM�ե��å����	*/
/*����������ߤ������ᡢHALT���DMAž���Ǥ��ʤ����꤫��pc_wait_flg�����ä���	*/
/*����������������pc_wait_flg��������Ƥξ�郎ɬ�פǤϤʤ����ᡢ		*/
/*��������stby_wait_flg�ξ��ˤ�����						*/
/*------------------------------------------------------------------------------*/
//	assign stby = (dec_halt | dec_stop) & ~stben & ~pc_wait_flg ;
	assign stby = (dec_halt | dec_stop) & ~stben & ~stby_wait_flg ;

// CPU������FLASH���򿮹��ޥ�������٤ο��档
// for EVA
//	assign flmask_pre = stby | waitfl | waitmod | waitexm | wait2ndsfr | waitint | waitdma ;
//	assign flmask_pre = stby | (waitfl | waitfl2 ) | waitmod | waitexm | wait2ndsfr | waitint | waitdma ;
	assign flmask_pre = stby | (waitfl | waitfl2 ) | waitmod | waitexm | wait2ndsfr | waitdflash | waitint | waitdma ;

//
	assign flmask = ~flmask_pre & cpustart ;

// ������Х����֤ȳ����������Ȥλ����Ȥʤ롣
// for EVA
//	assign cpuen_pre = flmask_pre ;
        assign cpuen_pre = flmask_pre | icewaitmem ;
//

// CPU���͡��֥뿮�档���ΤȤ�CPU����ߤ��롣
	assign cpuen = ~cpuen_pre & cpustart ;

// DMA�ѤΥ������ȿ��档
// for EVA
//	assign dmawait = waitexm | wait2ndsfr | waitfl | waitmod ;
//	assign dmawait = waitexm | wait2ndsfr | waitfl | waitmod | icewaitmem ;
	assign dmawait = waitexm | wait2ndsfr | waitdflash | waitfl | waitmod | icewaitmem ;
//

// OCD�ѤΥ������ȿ��档
	assign ocdwait = waitexm | wait2ndsfr | waitdflash ;

// RAM�ե��å����̿��ե��å�����(pc_wait_flg)��HALT/STOP������ʤ���
	assign hltst = ~pc_wait_flg & dec_halt ;
	assign stpst = ~pc_wait_flg & dec_stop ;

/*------------------------------------------------------------------------------*/
/* �꡼�ɥХ�									*/
/*------------------------------------------------------------------------------*/
/*   �ãУ���ӣƣҤΥ꡼�ɥХ��ȣң��ͤΥ꡼�ɥХ��Ȥ������¡�			*/
/*------------------------------------------------------------------------------*/

// CPU�������꡼�ɥХ���CPU��SFR�꡼�ɥХ��ȥ���꡼�ɥХ���OR��
	assign imdr = mdr | cpumdr ;

// for EVA
        assign cpumask = pselcpu & ((vpa == 4'h8) | (vpa == 4'h9) | (vpa == 4'ha) | (vpa == 4'hc) | (vpa == 4'hd)) ;
//

// for EVA
        assign SP_rd = (svmod & ~alt1) ? SP_sv : SP_usr ;
//

// CPU��SFR���쥸�����Х󥯤Υ꡼�ɥǡ�����
// for EVA
//	always @(pselcpu or cpurd or wdop or vpa or SP or PSW or CS or ES or MAA or
        always @(pselcpu or cpurd or wdop or vpa or SP_rd or PSW or CS or ES or MAA or
//
		 pselbcd or BCDADJ or slreg or rga or waitdma or
		 A_bank0 or X_bank0 or B_bank0 or C_bank0 or D_bank0 or E_bank0 or H_bank0 or L_bank0 or
		 A_bank1 or X_bank1 or B_bank1 or C_bank1 or D_bank1 or E_bank1 or H_bank1 or L_bank1 or
		 A_bank2 or X_bank2 or B_bank2 or C_bank2 or D_bank2 or E_bank2 or H_bank2 or L_bank2 or
		 A_bank3 or X_bank3 or B_bank3 or C_bank3 or D_bank3 or E_bank3 or H_bank3 or L_bank3 or
		RVEON ) begin
		if (waitdma) begin
			cpumdr = 16'h0000 ;
		end
		else if (pselcpu && cpurd) begin
			casex ({vpa,wdop})
// for EVA
//				({4'h8,1'b0}) : cpumdr = {8'h00,SP[6:0],1'b0} ;
//				({4'h8,1'b1}) : cpumdr = {SP,1'b0} ;
//				({4'h9,1'bx}) : cpumdr = {SP[14:7],8'h00} ;
                                ({4'h8,1'b0}) : cpumdr = {8'h00,SP_rd[6:0],1'b0} ;
                                ({4'h8,1'b1}) : cpumdr = {SP_rd,1'b0} ;
                                ({4'h9,1'bx}) : cpumdr = {SP_rd[14:7],8'h00} ;
//
				({4'ha,1'bx}) : cpumdr = {8'h00,PSW} ;
				({4'hc,1'b0}) : cpumdr = {12'h000,CS} ;
				({4'hc,1'b1}) : cpumdr = {4'h0,ES,4'h0,CS} ;
				({4'hd,1'bx}) : cpumdr = {4'h0,ES,8'h00} ;
				({4'he,1'bx}) : cpumdr = {15'b0,MAA} ;
				default : cpumdr = 16'h0000 ;
			endcase
		end
		else if (pselbcd && cpurd) begin
			casex ({vpa[0],wdop})
//				({1'b1,1'bx}) : cpumdr = {8'h00,8'h00} ;
//				({1'b0,1'b1}) : cpumdr = {8'h00,1'b0,BCDADJ[1],BCDADJ[1],1'b0,1'b0,BCDADJ[0],BCDADJ[0],1'b0} ;
				({1'b1,1'bx}) : cpumdr = {7'b0000_000,RVEON,8'h00} ;
				({1'b0,1'b0}) : cpumdr = {8'h00,1'b0,BCDADJ[1],BCDADJ[1],1'b0,1'b0,BCDADJ[0],BCDADJ[0],1'b0} ;
				({1'b0,1'b1}) : cpumdr = {7'b0000_000,RVEON,1'b0,BCDADJ[1],BCDADJ[1],1'b0,1'b0,BCDADJ[0],BCDADJ[0],1'b0} ;
				// cannot reach DEFAULT brunch
				// default : cpumdr = 16'h0000 ;
			endcase
		end
		else if (slreg && cpurd) begin
			casex ({rga,vpa,wdop})
				// ���إ쥸���� �Х󥯣�
				({1'b1,4'h9,1'bx}) : cpumdr = {A_bank0,8'h00  } ;
				({1'b1,4'h8,1'b0}) : cpumdr = {8'h00,  X_bank0} ;
				({1'b1,4'h8,1'b1}) : cpumdr = {A_bank0,X_bank0} ;
				// �£å쥸���� �Х󥯣�
				({1'b1,4'hb,1'bx}) : cpumdr = {B_bank0,8'h00  } ;
				({1'b1,4'ha,1'b0}) : cpumdr = {8'h00,  C_bank0} ;
				({1'b1,4'ha,1'b1}) : cpumdr = {B_bank0,C_bank0} ;
				// �ģť쥸���� �Х󥯣�
				({1'b1,4'hd,1'bx}) : cpumdr = {D_bank0,8'h00  } ;
				({1'b1,4'hc,1'b0}) : cpumdr = {8'h00,  E_bank0} ;
				({1'b1,4'hc,1'b1}) : cpumdr = {D_bank0,E_bank0} ;
				// �ȣ̥쥸���� �Х󥯣�
				({1'b1,4'hf,1'bx}) : cpumdr = {H_bank0,8'h00  } ;
				({1'b1,4'he,1'b0}) : cpumdr = {8'h00,  L_bank0} ;
				({1'b1,4'he,1'b1}) : cpumdr = {H_bank0,L_bank0} ;
				// ���إ쥸���� �Х󥯣�
				({1'b1,4'h1,1'bx}) : cpumdr = {A_bank1,8'h00  } ;
				({1'b1,4'h0,1'b0}) : cpumdr = {8'h00,  X_bank1} ;
				({1'b1,4'h0,1'b1}) : cpumdr = {A_bank1,X_bank1} ;
				// �£å쥸���� �Х󥯣�
				({1'b1,4'h3,1'bx}) : cpumdr = {B_bank1,8'h00  } ;
				({1'b1,4'h2,1'b0}) : cpumdr = {8'h00,  C_bank1} ;
				({1'b1,4'h2,1'b1}) : cpumdr = {B_bank1,C_bank1} ;
				// �ģť쥸���� �Х󥯣�
				({1'b1,4'h5,1'bx}) : cpumdr = {D_bank1,8'h00  } ;
				({1'b1,4'h4,1'b0}) : cpumdr = {8'h00,  E_bank1} ;
				({1'b1,4'h4,1'b1}) : cpumdr = {D_bank1,E_bank1} ;
				// �ȣ̥쥸���� �Х󥯣�
				({1'b1,4'h7,1'bx}) : cpumdr = {H_bank1,8'h00  } ;
				({1'b1,4'h6,1'b0}) : cpumdr = {8'h00,  L_bank1} ;
				({1'b1,4'h6,1'b1}) : cpumdr = {H_bank1,L_bank1} ;
				// ���إ쥸���� �Х󥯣�
				({1'b0,4'h9,1'bx}) : cpumdr = {A_bank2,8'h00  } ;
				({1'b0,4'h8,1'b0}) : cpumdr = {8'h00,  X_bank2} ;
				({1'b0,4'h8,1'b1}) : cpumdr = {A_bank2,X_bank2} ;
				// �£å쥸���� �Х󥯣�
				({1'b0,4'hb,1'bx}) : cpumdr = {B_bank2,8'h00  } ;
				({1'b0,4'ha,1'b0}) : cpumdr = {8'h00,  C_bank2} ;
				({1'b0,4'ha,1'b1}) : cpumdr = {B_bank2,C_bank2} ;
				// �ģť쥸���� �Х󥯣�
				({1'b0,4'hd,1'bx}) : cpumdr = {D_bank2,8'h00  } ;
				({1'b0,4'hc,1'b0}) : cpumdr = {8'h00,  E_bank2} ;
				({1'b0,4'hc,1'b1}) : cpumdr = {D_bank2,E_bank2} ;
				// �ȣ̥쥸���� �Х󥯣�
				({1'b0,4'hf,1'bx}) : cpumdr = {H_bank2,8'h00  } ;
				({1'b0,4'he,1'b0}) : cpumdr = {8'h00,  L_bank2} ;
				({1'b0,4'he,1'b1}) : cpumdr = {H_bank2,L_bank2} ;
				// ���إ쥸���� �Х󥯣�
				({1'b0,4'h1,1'bx}) : cpumdr = {A_bank3,8'h00  } ;
				({1'b0,4'h0,1'b0}) : cpumdr = {8'h00,  X_bank3} ;
				({1'b0,4'h0,1'b1}) : cpumdr = {A_bank3,X_bank3} ;
				// �£å쥸���� �Х󥯣�
				({1'b0,4'h3,1'bx}) : cpumdr = {B_bank3,8'h00  } ;
				({1'b0,4'h2,1'b0}) : cpumdr = {8'h00,  C_bank3} ;
				({1'b0,4'h2,1'b1}) : cpumdr = {B_bank3,C_bank3} ;
				// �ģť쥸���� �Х󥯣�
				({1'b0,4'h5,1'bx}) : cpumdr = {D_bank3,8'h00  } ;
				({1'b0,4'h4,1'b0}) : cpumdr = {8'h00,  E_bank3} ;
				({1'b0,4'h4,1'b1}) : cpumdr = {D_bank3,E_bank3} ;
				// �ȣ̥쥸���� �Х󥯣�
				({1'b0,4'h7,1'bx}) : cpumdr = {H_bank3,8'h00  } ;
				({1'b0,4'h6,1'b0}) : cpumdr = {8'h00,  L_bank3} ;
				({1'b0,4'h6,1'b1}) : cpumdr = {H_bank3,L_bank3} ;
				// cannot reach DEFAULT brunch
				// default : cpumdr = 16'h0000 ;
			endcase
		end
		else cpumdr = 16'h0000 ;
	end

endmodule

/************************************************************************/
/* Module Name : QLK0RCPUEVA0V3_DEC                                        */
/* Author      : K.Kawai                                                */
/* Rev, Date   : 1.0 2006/1/13 11:41:29 generated by make_superk0.c.    */
/************************************************************************/

module QLK0RCPUEVA0V3_DEC(
        ID_stage1, /* ID Code address stage 15-8bit */
        ID_stage0, /* ID Code address stage 7-0bit */
        stage_adr,         /* Address stage machine cycle */
        rstvec,             /* RESET Vector */
        ivack,             /* Interrupt Vector ACK */
        skpack,             /* Skip ACK */
        dec_alu_input10,   /* ALU input1[7:0] */
        dec_alu_input20,   /* ALU input2[7:0] */
        dec_alu_add,    
        dec_alu_sub,    
        dec_alu_and,    
        dec_alu_or,    
        dec_alu_exor,    
        dec_alu_andbit,    
        dec_alu_orbit,    
        dec_alu_exorbit,    
        dec_alu_ror,    
        dec_alu_rol,    
        dec_alu_shr,    
        dec_alu_shl,    
        dec_alu_sar,    
        dec_alu_mulu,    
        dec_alu_carry,    
	dec_alu_transout,  /* trans instruction MOV,XCH,MOVW,XCHW */
	dec_alu_transin,   /* trans instruction MOV,XCH,MOVW,XCHW */
	dec_alu_bitsh,  /* bit,shift instruction ROR, SHR, MOV1, AND1, etc... */
	dec_alu_biten,	/* biten instruction */
        dec_word_access,   /* Word access */
        dec_xch_byte,      /* XCH resister direct input byte */
        dec_xchw_bc,       /* XCHW resister direct input AX<-BC */
        dec_xchw_de,       /* XCHW resister direct input AX<-DE */
        dec_xchw_hl,       /* XCHW resister direct input AX<-HL */
        dec_SP_enable,
        dec_A_enable,
        dec_X_enable,
        dec_B_enable,
        dec_C_enable,
        dec_D_enable,
        dec_E_enable,
        dec_H_enable,
        dec_L_enable,
        dec_ES_enable,
        dec_Z_enable,
        dec_CY_enable,
        dec_AC_enable,
        dec_IE_enable,
        dec_ISP_enable,
        dec_RBS_enable,
        dec_NMIS_enable,
        dec_buf0_enable,
        dec_buf1_enable,
        dec_buf2_enable,
        dec_cpuwr_enable,
        dec_cpurd_enable,
        dec_ma_enable,
        dec_ma_data_sp,
        dec_ma_data_saddr_op1,
        dec_ma_data_saddr_op2,
        dec_ma_data_sfr_op1,
        dec_ma_data_sfr_op2,
        dec_ma_data_op12,
        dec_ma_data_op23,
        dec_ma_data_HL,
        dec_ma_data_HLop1,
        dec_ma_data_HLop2,
        dec_ma_data_HLB,
        dec_ma_data_HLC,
        dec_ma_data_DE,
        dec_ma_data_DEop1,
        dec_ma_data_DEop2,
        dec_ma_data_SPop1,
        dec_ma_data_BCop12,
        dec_ma_data_Bop12,
        dec_ma_data_Cop12,
        dec_sp_set_enable,
        dec_sp_inc,
        dec_sp_dec,
        dec_pc_inc1,
        dec_pc_inc2,
        dec_pc_inc3,
        dec_pc_inc4,
        dec_clear_stage,
        dec_pc_set_enable,
        dec_pc_set_op01,
        dec_pc_set_op12,
        dec_pc_set_op123,
        dec_pc_set_AX,
        dec_pc_set_BC,
        dec_pc_set_DE,
        dec_pc_set_HL,
        dec_pc_set_pc1,
        dec_pc_set_pc2,
        dec_pc_set_pc3,
        dec_pc_set_pc12,
        dec_pc_set_calt,
        dec_pc_set_vec,
        dec_pc_set_brk,
        dec_pc_set_dbg,
        dec_pc_set_ret,
        dec_stage_cut_brtf,
        dec_stage_cut_ifbr,
        dec_ifbr_not,
        dec_ifbr_zero,
        dec_ifbr_ht,
        dec_mem_stage_op2,
        dec_mem_stage_op3,
        dec_mem_stage_op23,
        dec_set_buf_retadr,
        dec_set_buf_intr,
        dec_skc,
        dec_sknc,
        dec_skz,
        dec_sknz,
        dec_skh,
        dec_sknh,
        dec_prefix,
        dec_halt,
        dec_stop,
        dec_movs,
        dec_cmps,
// for EVA
        dec_alt1,
        dec_alt2,
//
        baseck, resb,scanmode,cpuen);
    input [7:0] ID_stage1, ID_stage0;
    input [1:0] stage_adr;
    input       rstvec;
    input       ivack;
    input       skpack;
    input       baseck, resb,scanmode,cpuen;

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����������ɥ쥹���ơ����Υǥ��������Ϥϡ��ǥ������ΥХ��Ĥ������Τޤ޽��Ϥ�	*/
/*����������롣���ΥХ��Ĥ��ˤ����ή��︺����٤ˡ��ǥ��������Ϥ�Ƭ��	*/
/*���������ޥ��������ϩ���������롣�����������ԡ��ɥͥå��Ȥʤ뤿��		*/
/*��������(�ǥ��������Ϣ�SLFLASH)��AMPH=1�λ��ϥѥ������롣			*/
/*------------------------------------------------------------------------------*/
/* Ver3.0 �ǥ��쥤�ˤ��ҥ��ɻ߲�ϩ���к���ľ��(CPUv1.5���������᤹)		*/
/*------------------------------------------------------------------------------*/

//    wire decout_mask, decout_mask_dly;
//    QLK0RCPUEVA0V3_DEC_DLY dec_delay (.out(decout_mask_dly), .in(decout_mask_reg));
//    assign decout_mask = decout_mask_reg ^ (decout_mask_dly & ~scanmode);

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*����INC,DEC,INCW,DECW,ADD,ADDC,SUB,SUBC,AND,OR,XOR�Υ��ꥢ�������黻��	*/
/*������������å��ܤ��飱����å��ܤ��ѹ���					*/
/*�����ӥå����̿�ᡢBT,BF,BTCLR�����̺����dec_alu_bitsh�ذ�ư		*/
/*����ONE̿������̺����dec_alu_transout�ذ�ư					*/
/*����MULU̿�������dec_alu_mulu�ذ�ư					*/
/*------------------------------------------------------------------------------*/

    output [3:0] dec_alu_input10;
    reg    [3:0] dec_alu_input10, dec_alu_input10_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_alu_input10_adrstage = 4'h0;
        end else begin
            if(ID_stage0 == 8'h61) begin
                casex ({ID_stage1,stage_adr})  
                    {8'h08,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADD,A,X */
                    {8'h0a,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADD,A,C */
                    {8'h0b,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADD,A,B */
                    {8'h0c,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADD,A,E */
                    {8'h0d,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADD,A,D */
                    {8'h0e,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADD,A,L */
                    {8'h0f,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADD,A,H */
                    {8'h00,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* ADD,X,A */
                    {8'h01,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADD,A,A */
                    {8'h02,2'bxx} : dec_alu_input10_adrstage = 4'h6;  /* ADD,C,A */
                    {8'h03,2'bxx} : dec_alu_input10_adrstage = 4'h5;  /* ADD,B,A */
                    {8'h04,2'bxx} : dec_alu_input10_adrstage = 4'h8;  /* ADD,E,A */
                    {8'h05,2'bxx} : dec_alu_input10_adrstage = 4'h7;  /* ADD,D,A */
                    {8'h06,2'bxx} : dec_alu_input10_adrstage = 4'ha;  /* ADD,L,A */
                    {8'h07,2'bxx} : dec_alu_input10_adrstage = 4'h9;  /* ADD,H,A */
                    {8'h80,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADD,A,[HL+B] */
                    {8'h82,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADD,A,[HL+C] */
                    {8'h18,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADDC,A,X */
                    {8'h1a,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADDC,A,C */
                    {8'h1b,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADDC,A,B */
                    {8'h1c,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADDC,A,E */
                    {8'h1d,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADDC,A,D */
                    {8'h1e,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADDC,A,L */
                    {8'h1f,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADDC,A,H */
                    {8'h10,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* ADDC,X,A */
                    {8'h11,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADDC,A,A */
                    {8'h12,2'bxx} : dec_alu_input10_adrstage = 4'h6;  /* ADDC,C,A */
                    {8'h13,2'bxx} : dec_alu_input10_adrstage = 4'h5;  /* ADDC,B,A */
                    {8'h14,2'bxx} : dec_alu_input10_adrstage = 4'h8;  /* ADDC,E,A */
                    {8'h15,2'bxx} : dec_alu_input10_adrstage = 4'h7;  /* ADDC,D,A */
                    {8'h16,2'bxx} : dec_alu_input10_adrstage = 4'ha;  /* ADDC,L,A */
                    {8'h17,2'bxx} : dec_alu_input10_adrstage = 4'h9;  /* ADDC,H,A */
                    {8'h90,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADDC,A,[HL+B] */
                    {8'h92,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADDC,A,[HL+C] */
                    {8'h28,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUB,A,X */
                    {8'h2a,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUB,A,C */
                    {8'h2b,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUB,A,B */
                    {8'h2c,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUB,A,E */
                    {8'h2d,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUB,A,D */
                    {8'h2e,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUB,A,L */
                    {8'h2f,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUB,A,H */
                    {8'h20,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* SUB,X,A */
                    {8'h21,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUB,A,A */
                    {8'h22,2'bxx} : dec_alu_input10_adrstage = 4'h6;  /* SUB,C,A */
                    {8'h23,2'bxx} : dec_alu_input10_adrstage = 4'h5;  /* SUB,B,A */
                    {8'h24,2'bxx} : dec_alu_input10_adrstage = 4'h8;  /* SUB,E,A */
                    {8'h25,2'bxx} : dec_alu_input10_adrstage = 4'h7;  /* SUB,D,A */
                    {8'h26,2'bxx} : dec_alu_input10_adrstage = 4'ha;  /* SUB,L,A */
                    {8'h27,2'bxx} : dec_alu_input10_adrstage = 4'h9;  /* SUB,H,A */
                    {8'ha0,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUB,A,[HL+B] */
                    {8'ha2,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUB,A,[HL+C] */
                    {8'h38,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUBC,A,X */
                    {8'h3a,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUBC,A,C */
                    {8'h3b,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUBC,A,B */
                    {8'h3c,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUBC,A,E */
                    {8'h3d,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUBC,A,D */
                    {8'h3e,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUBC,A,L */
                    {8'h3f,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUBC,A,H */
                    {8'h30,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* SUBC,X,A */
                    {8'h31,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUBC,A,A */
                    {8'h32,2'bxx} : dec_alu_input10_adrstage = 4'h6;  /* SUBC,C,A */
                    {8'h33,2'bxx} : dec_alu_input10_adrstage = 4'h5;  /* SUBC,B,A */
                    {8'h34,2'bxx} : dec_alu_input10_adrstage = 4'h8;  /* SUBC,E,A */
                    {8'h35,2'bxx} : dec_alu_input10_adrstage = 4'h7;  /* SUBC,D,A */
                    {8'h36,2'bxx} : dec_alu_input10_adrstage = 4'ha;  /* SUBC,L,A */
                    {8'h37,2'bxx} : dec_alu_input10_adrstage = 4'h9;  /* SUBC,H,A */
                    {8'hb0,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUBC,A,[HL+B] */
                    {8'hb2,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUBC,A,[HL+C] */
                    {8'h58,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* AND,A,X */
                    {8'h5a,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* AND,A,C */
                    {8'h5b,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* AND,A,B */
                    {8'h5c,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* AND,A,E */
                    {8'h5d,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* AND,A,D */
                    {8'h5e,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* AND,A,L */
                    {8'h5f,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* AND,A,H */
                    {8'h50,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* AND,X,A */
                    {8'h51,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* AND,A,A */
                    {8'h52,2'bxx} : dec_alu_input10_adrstage = 4'h6;  /* AND,C,A */
                    {8'h53,2'bxx} : dec_alu_input10_adrstage = 4'h5;  /* AND,B,A */
                    {8'h54,2'bxx} : dec_alu_input10_adrstage = 4'h8;  /* AND,E,A */
                    {8'h55,2'bxx} : dec_alu_input10_adrstage = 4'h7;  /* AND,D,A */
                    {8'h56,2'bxx} : dec_alu_input10_adrstage = 4'ha;  /* AND,L,A */
                    {8'h57,2'bxx} : dec_alu_input10_adrstage = 4'h9;  /* AND,H,A */
                    {8'hd0,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* AND,A,[HL+B] */
                    {8'hd2,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* AND,A,[HL+C] */
                    {8'h68,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* OR,A,X */
                    {8'h6a,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* OR,A,C */
                    {8'h6b,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* OR,A,B */
                    {8'h6c,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* OR,A,E */
                    {8'h6d,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* OR,A,D */
                    {8'h6e,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* OR,A,L */
                    {8'h6f,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* OR,A,H */
                    {8'h60,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* OR,X,A */
                    {8'h61,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* OR,A,A */
                    {8'h62,2'bxx} : dec_alu_input10_adrstage = 4'h6;  /* OR,C,A */
                    {8'h63,2'bxx} : dec_alu_input10_adrstage = 4'h5;  /* OR,B,A */
                    {8'h64,2'bxx} : dec_alu_input10_adrstage = 4'h8;  /* OR,E,A */
                    {8'h65,2'bxx} : dec_alu_input10_adrstage = 4'h7;  /* OR,D,A */
                    {8'h66,2'bxx} : dec_alu_input10_adrstage = 4'ha;  /* OR,L,A */
                    {8'h67,2'bxx} : dec_alu_input10_adrstage = 4'h9;  /* OR,H,A */
                    {8'he0,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* OR,A,[HL+B] */
                    {8'he2,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* OR,A,[HL+C] */
                    {8'h78,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* XOR,A,X */
                    {8'h7a,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* XOR,A,C */
                    {8'h7b,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* XOR,A,B */
                    {8'h7c,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* XOR,A,E */
                    {8'h7d,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* XOR,A,D */
                    {8'h7e,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* XOR,A,L */
                    {8'h7f,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* XOR,A,H */
                    {8'h70,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* XOR,X,A */
                    {8'h71,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* XOR,A,A */
                    {8'h72,2'bxx} : dec_alu_input10_adrstage = 4'h6;  /* XOR,C,A */
                    {8'h73,2'bxx} : dec_alu_input10_adrstage = 4'h5;  /* XOR,B,A */
                    {8'h74,2'bxx} : dec_alu_input10_adrstage = 4'h8;  /* XOR,E,A */
                    {8'h75,2'bxx} : dec_alu_input10_adrstage = 4'h7;  /* XOR,D,A */
                    {8'h76,2'bxx} : dec_alu_input10_adrstage = 4'ha;  /* XOR,L,A */
                    {8'h77,2'bxx} : dec_alu_input10_adrstage = 4'h9;  /* XOR,H,A */
                    {8'hf0,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* XOR,A,[HL+B] */
                    {8'hf2,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* XOR,A,[HL+C] */
                    {8'h48,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* CMP,A,X */
                    {8'h4a,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* CMP,A,C */
                    {8'h4b,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* CMP,A,B */
                    {8'h4c,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* CMP,A,E */
                    {8'h4d,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* CMP,A,D */
                    {8'h4e,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* CMP,A,L */
                    {8'h4f,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* CMP,A,H */
                    {8'h40,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* CMP,X,A */
                    {8'h41,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* CMP,A,A */
                    {8'h42,2'bxx} : dec_alu_input10_adrstage = 4'h6;  /* CMP,C,A */
                    {8'h43,2'bxx} : dec_alu_input10_adrstage = 4'h5;  /* CMP,B,A */
                    {8'h44,2'bxx} : dec_alu_input10_adrstage = 4'h8;  /* CMP,E,A */
                    {8'h45,2'bxx} : dec_alu_input10_adrstage = 4'h7;  /* CMP,D,A */
                    {8'h46,2'bxx} : dec_alu_input10_adrstage = 4'ha;  /* CMP,L,A */
                    {8'h47,2'bxx} : dec_alu_input10_adrstage = 4'h9;  /* CMP,H,A */
                    {8'hc0,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* CMP,A,[HL+B] */
                    {8'hc2,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* CMP,A,[HL+C] */
                    {8'hde,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* CMPS,X,[HL+byte] */
                    {8'h09,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* ADDW,AX,[HL+byte] */
                    {8'h29,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* SUBW,AX,[HL+byte] */
                    {8'h49,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* CMPW,AX,[HL+byte] */
                    {8'h59,2'bx0} : dec_alu_input10_adrstage = 4'hb;  /* INC,,[HL+byte] */
                    {8'h69,2'bx0} : dec_alu_input10_adrstage = 4'hb;  /* DEC,,[HL+byte] */
                    {8'h79,2'bx0} : dec_alu_input10_adrstage = 4'hb;  /* INCW,,[HL+byte] */
                    {8'h89,2'bx0} : dec_alu_input10_adrstage = 4'hb;  /* DECW,,[HL+byte] */
                    {8'h19,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADDC,A,A */
                    {8'h39,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUBC,A,A */
                    {8'hd1,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* AND,A,[HL+B] */
                    {8'he1,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* OR,A,[HL+B] */
                    {8'hf1,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* XOR,A,[HL+B] */
                    {8'h83,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADD,A,[HL+C] */
                    {8'h93,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADDC,A,[HL+C] */
                    {8'ha3,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUB,A,[HL+C] */
                    {8'hb3,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUBC,A,[HL+C] */
                    default : dec_alu_input10_adrstage = 4'h0;
                endcase
            end else if(ID_stage0 == 8'h71) begin
                    dec_alu_input10_adrstage = 4'h0;
            end else if(ID_stage0 == 8'h31) begin
                    dec_alu_input10_adrstage = 4'h0;
            end else begin
                casex ({ID_stage0,stage_adr})  
                    {8'h0c,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADD,A,#byte */
                    {8'h0a,2'bx0} : dec_alu_input10_adrstage = 4'he;  /* ADD,saddr,#byte */
                    {8'h0b,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADD,A,saddr */
                    {8'h0f,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADD,A,!addr16 */
                    {8'h0d,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADD,A,[HL] */
                    {8'h0e,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADD,A,[HL+byte] */
                    {8'h1c,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADDC,A,#byte */
                    {8'h1a,2'bx0} : dec_alu_input10_adrstage = 4'he;  /* ADDC,saddr,#byte */
                    {8'h1b,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADDC,A,saddr */
                    {8'h1f,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADDC,A,!addr16 */
                    {8'h1d,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADDC,A,[HL] */
                    {8'h1e,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* ADDC,A,[HL+byte] */
                    {8'h2c,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUB,A,#byte */
                    {8'h2a,2'bx0} : dec_alu_input10_adrstage = 4'he;  /* SUB,saddr,#byte */
                    {8'h2b,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUB,A,saddr */
                    {8'h2f,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUB,A,!addr16 */
                    {8'h2d,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUB,A,[HL] */
                    {8'h2e,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUB,A,[HL+byte] */
                    {8'h3c,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUBC,A,#byte */
                    {8'h3a,2'bx0} : dec_alu_input10_adrstage = 4'he;  /* SUBC,saddr,#byte */
                    {8'h3b,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUBC,A,saddr */
                    {8'h3f,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUBC,A,!addr16 */
                    {8'h3d,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUBC,A,[HL] */
                    {8'h3e,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* SUBC,A,[HL+byte] */
                    {8'h5c,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* AND,A,#byte */
                    {8'h5a,2'bx0} : dec_alu_input10_adrstage = 4'he;  /* AND,saddr,#byte */
                    {8'h5b,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* AND,A,saddr */
                    {8'h5f,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* AND,A,!addr16 */
                    {8'h5d,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* AND,A,[HL] */
                    {8'h5e,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* AND,A,[HL+byte] */
                    {8'h6c,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* OR,A,#byte */
                    {8'h6a,2'bx0} : dec_alu_input10_adrstage = 4'he;  /* OR,saddr,#byte */
                    {8'h6b,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* OR,A,saddr */
                    {8'h6f,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* OR,A,!addr16 */
                    {8'h6d,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* OR,A,[HL] */
                    {8'h6e,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* OR,A,[HL+byte] */
                    {8'h7c,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* XOR,A,#byte */
                    {8'h7a,2'bx0} : dec_alu_input10_adrstage = 4'he;  /* XOR,saddr,#byte */
                    {8'h7b,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* XOR,A,saddr */
                    {8'h7f,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* XOR,A,!addr16 */
                    {8'h7d,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* XOR,A,[HL] */
                    {8'h7e,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* XOR,A,[HL+byte] */
                    {8'h4c,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* CMP,A,#byte */
                    {8'h4a,2'bxx} : dec_alu_input10_adrstage = 4'he;  /* CMP,saddr,#byte */
                    {8'h40,2'bxx} : dec_alu_input10_adrstage = 4'he;  /* CMP,!addr16,#byte */
                    {8'h4b,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* CMP,A,saddr */
                    {8'h4f,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* CMP,A,!addr16 */
                    {8'h4d,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* CMP,A,[HL] */
                    {8'h4e,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* CMP,A,[HL+byte] */
                    {8'hd1,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* CMP0,,A */
                    {8'hd0,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* CMP0,,X */
                    {8'hd3,2'bxx} : dec_alu_input10_adrstage = 4'h5;  /* CMP0,,B */
                    {8'hd2,2'bxx} : dec_alu_input10_adrstage = 4'h6;  /* CMP0,,C */
                    {8'hd4,2'bxx} : dec_alu_input10_adrstage = 4'he;  /* CMP0,,saddr */
                    {8'hd5,2'bxx} : dec_alu_input10_adrstage = 4'he;  /* CMP0,,!addr16 */
                    {8'h04,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* ADDW,AX,#word */
                    {8'h01,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* ADDW,AX,AX */
                    {8'h03,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* ADDW,AX,BC */
                    {8'h05,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* ADDW,AX,DE */
                    {8'h07,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* ADDW,AX,HL */
                    {8'h06,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* ADDW,AX,saddrp */
                    {8'h02,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* ADDW,AX,!addr16 */
                    {8'h24,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* SUBW,AX,#word */
                    {8'h21,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* SUBW,AX,AX */
                    {8'h23,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* SUBW,AX,BC */
                    {8'h25,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* SUBW,AX,DE */
                    {8'h27,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* SUBW,AX,HL */
                    {8'h26,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* SUBW,AX,saddrp */
                    {8'h22,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* SUBW,AX,!addr16 */
                    {8'h44,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* CMPW,AX,#word */
                    {8'h43,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* CMPW,AX,BC */
                    {8'h45,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* CMPW,AX,DE */
                    {8'h47,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* CMPW,AX,HL */
                    {8'h46,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* CMPW,AX,saddrp */
                    {8'h42,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* CMPW,AX,!addr16 */
                    {8'h80,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* INC,,X */
                    {8'h81,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* INC,,A */
                    {8'h82,2'bxx} : dec_alu_input10_adrstage = 4'h6;  /* INC,,C */
                    {8'h83,2'bxx} : dec_alu_input10_adrstage = 4'h5;  /* INC,,B */
                    {8'h84,2'bxx} : dec_alu_input10_adrstage = 4'h8;  /* INC,,E */
                    {8'h85,2'bxx} : dec_alu_input10_adrstage = 4'h7;  /* INC,,D */
                    {8'h86,2'bxx} : dec_alu_input10_adrstage = 4'ha;  /* INC,,L */
                    {8'h87,2'bxx} : dec_alu_input10_adrstage = 4'h9;  /* INC,,H */
                    {8'ha4,2'bx0} : dec_alu_input10_adrstage = 4'he;  /* INC,,saddr */
                    {8'ha0,2'bx0} : dec_alu_input10_adrstage = 4'he;  /* INC,,!addr16 */
                    {8'h90,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* DEC,,X */
                    {8'h91,2'bxx} : dec_alu_input10_adrstage = 4'h3;  /* DEC,,A */
                    {8'h92,2'bxx} : dec_alu_input10_adrstage = 4'h6;  /* DEC,,C */
                    {8'h93,2'bxx} : dec_alu_input10_adrstage = 4'h5;  /* DEC,,B */
                    {8'h94,2'bxx} : dec_alu_input10_adrstage = 4'h8;  /* DEC,,E */
                    {8'h95,2'bxx} : dec_alu_input10_adrstage = 4'h7;  /* DEC,,D */
                    {8'h96,2'bxx} : dec_alu_input10_adrstage = 4'ha;  /* DEC,,L */
                    {8'h97,2'bxx} : dec_alu_input10_adrstage = 4'h9;  /* DEC,,H */
                    {8'hb4,2'bx0} : dec_alu_input10_adrstage = 4'he;  /* DEC,,saddr */
                    {8'hb0,2'bx0} : dec_alu_input10_adrstage = 4'he;  /* DEC,,!addr16 */
                    {8'ha1,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* INCW,,AX */
                    {8'ha3,2'bxx} : dec_alu_input10_adrstage = 4'h6;  /* INCW,,BC */
                    {8'ha5,2'bxx} : dec_alu_input10_adrstage = 4'h8;  /* INCW,,DE */
                    {8'ha7,2'bxx} : dec_alu_input10_adrstage = 4'ha;  /* INCW,,HL */
                    {8'ha6,2'bx0} : dec_alu_input10_adrstage = 4'hb;  /* INCW,,saddrp */
                    {8'ha2,2'bx0} : dec_alu_input10_adrstage = 4'hb;  /* INCW,,!addr16 */
                    {8'hb1,2'bxx} : dec_alu_input10_adrstage = 4'h4;  /* DECW,,AX */
                    {8'hb3,2'bxx} : dec_alu_input10_adrstage = 4'h6;  /* DECW,,BC */
                    {8'hb5,2'bxx} : dec_alu_input10_adrstage = 4'h8;  /* DECW,,DE */
                    {8'hb7,2'bxx} : dec_alu_input10_adrstage = 4'ha;  /* DECW,,HL */
                    {8'hb6,2'bx0} : dec_alu_input10_adrstage = 4'he;  /* DECW,,saddrp */
                    {8'hb2,2'bx0} : dec_alu_input10_adrstage = 4'he;  /* DECW,,!addr16 */
                    {8'h10,2'bxx} : dec_alu_input10_adrstage = 4'hd;  /* ADDW,SP,#byte */
                    {8'h20,2'bxx} : dec_alu_input10_adrstage = 4'hd;  /* SUBW,SP,#byte */
                    default : dec_alu_input10_adrstage = 4'h0;
                endcase
            end
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_alu_input10 <= 4'h0;
        else if(cpuen) dec_alu_input10 <= dec_alu_input10_adrstage;
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*����MOV,MOVS,MOVW,XCH,XCHW̿������̺����dec_alu_transin,			*/
/*							dec_alu_trans_out�ذ�ư	*/
/*    ROR,ROL,RORC,ROLC,ROLWC�����̺����dec_alu_bitsh�ذ�ư			*/
/*����CALL,CALLT,BRK,SOFT,PUSH�����̺����dec_alu_transout�ذ�ư		*/
/*�����ӥå����̿�ᡢBT,BF,BTCLR�����̺����dec_alu_bitsh�ذ�ư		*/
/*����SHR,SHRW,SHL,SHLW,SAR,SARW�����̺����dec_alu_bitsh�ذ�ư			*/
/*����MULU̿�������dec_alu_mulu�ذ�ư					*/
/*������郎���ä����ᡢ5bit��4bit���ѹ�					*/
/*------------------------------------------------------------------------------*/

    output [3:0] dec_alu_input20;
    reg    [3:0] dec_alu_input20, dec_alu_input20_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_alu_input20_adrstage = 4'h0;
        end else begin
            if(ID_stage0 == 8'h61) begin
                casex ({ID_stage1,stage_adr})  
                    {8'h08,2'bxx} : dec_alu_input20_adrstage = 4'h3;  /* ADD,A,X */
                    {8'h0a,2'bxx} : dec_alu_input20_adrstage = 4'h5;  /* ADD,A,C */
                    {8'h0b,2'bxx} : dec_alu_input20_adrstage = 4'h4;  /* ADD,A,B */
                    {8'h0c,2'bxx} : dec_alu_input20_adrstage = 4'h7;  /* ADD,A,E */
                    {8'h0d,2'bxx} : dec_alu_input20_adrstage = 4'h6;  /* ADD,A,D */
                    {8'h0e,2'bxx} : dec_alu_input20_adrstage = 4'h9;  /* ADD,A,L */
                    {8'h0f,2'bxx} : dec_alu_input20_adrstage = 4'h8;  /* ADD,A,H */
                    {8'h00,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* ADD,X,A */
                    {8'h01,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* ADD,A,A */
                    {8'h02,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* ADD,C,A */
                    {8'h03,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* ADD,B,A */
                    {8'h04,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* ADD,E,A */
                    {8'h05,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* ADD,D,A */
                    {8'h06,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* ADD,L,A */
                    {8'h07,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* ADD,H,A */
                    {8'h80,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* ADD,A,[HL+B] */
                    {8'h82,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* ADD,A,[HL+C] */
                    {8'h18,2'bxx} : dec_alu_input20_adrstage = 4'h3;  /* ADDC,A,X */
                    {8'h1a,2'bxx} : dec_alu_input20_adrstage = 4'h5;  /* ADDC,A,C */
                    {8'h1b,2'bxx} : dec_alu_input20_adrstage = 4'h4;  /* ADDC,A,B */
                    {8'h1c,2'bxx} : dec_alu_input20_adrstage = 4'h7;  /* ADDC,A,E */
                    {8'h1d,2'bxx} : dec_alu_input20_adrstage = 4'h6;  /* ADDC,A,D */
                    {8'h1e,2'bxx} : dec_alu_input20_adrstage = 4'h9;  /* ADDC,A,L */
                    {8'h1f,2'bxx} : dec_alu_input20_adrstage = 4'h8;  /* ADDC,A,H */
                    {8'h10,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* ADDC,X,A */
                    {8'h11,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* ADDC,A,A */
                    {8'h12,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* ADDC,C,A */
                    {8'h13,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* ADDC,B,A */
                    {8'h14,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* ADDC,E,A */
                    {8'h15,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* ADDC,D,A */
                    {8'h16,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* ADDC,L,A */
                    {8'h17,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* ADDC,H,A */
                    {8'h90,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* ADDC,A,[HL+B] */
                    {8'h92,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* ADDC,A,[HL+C] */
                    {8'h28,2'bxx} : dec_alu_input20_adrstage = 4'h3;  /* SUB,A,X */
                    {8'h2a,2'bxx} : dec_alu_input20_adrstage = 4'h5;  /* SUB,A,C */
                    {8'h2b,2'bxx} : dec_alu_input20_adrstage = 4'h4;  /* SUB,A,B */
                    {8'h2c,2'bxx} : dec_alu_input20_adrstage = 4'h7;  /* SUB,A,E */
                    {8'h2d,2'bxx} : dec_alu_input20_adrstage = 4'h6;  /* SUB,A,D */
                    {8'h2e,2'bxx} : dec_alu_input20_adrstage = 4'h9;  /* SUB,A,L */
                    {8'h2f,2'bxx} : dec_alu_input20_adrstage = 4'h8;  /* SUB,A,H */
                    {8'h20,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* SUB,X,A */
                    {8'h21,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* SUB,A,A */
                    {8'h22,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* SUB,C,A */
                    {8'h23,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* SUB,B,A */
                    {8'h24,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* SUB,E,A */
                    {8'h25,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* SUB,D,A */
                    {8'h26,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* SUB,L,A */
                    {8'h27,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* SUB,H,A */
                    {8'ha0,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* SUB,A,[HL+B] */
                    {8'ha2,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* SUB,A,[HL+C] */
                    {8'h38,2'bxx} : dec_alu_input20_adrstage = 4'h3;  /* SUBC,A,X */
                    {8'h3a,2'bxx} : dec_alu_input20_adrstage = 4'h5;  /* SUBC,A,C */
                    {8'h3b,2'bxx} : dec_alu_input20_adrstage = 4'h4;  /* SUBC,A,B */
                    {8'h3c,2'bxx} : dec_alu_input20_adrstage = 4'h7;  /* SUBC,A,E */
                    {8'h3d,2'bxx} : dec_alu_input20_adrstage = 4'h6;  /* SUBC,A,D */
                    {8'h3e,2'bxx} : dec_alu_input20_adrstage = 4'h9;  /* SUBC,A,L */
                    {8'h3f,2'bxx} : dec_alu_input20_adrstage = 4'h8;  /* SUBC,A,H */
                    {8'h30,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* SUBC,X,A */
                    {8'h31,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* SUBC,A,A */
                    {8'h32,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* SUBC,C,A */
                    {8'h33,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* SUBC,B,A */
                    {8'h34,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* SUBC,E,A */
                    {8'h35,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* SUBC,D,A */
                    {8'h36,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* SUBC,L,A */
                    {8'h37,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* SUBC,H,A */
                    {8'hb0,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* SUBC,A,[HL+B] */
                    {8'hb2,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* SUBC,A,[HL+C] */
                    {8'h58,2'bxx} : dec_alu_input20_adrstage = 4'h3;  /* AND,A,X */
                    {8'h5a,2'bxx} : dec_alu_input20_adrstage = 4'h5;  /* AND,A,C */
                    {8'h5b,2'bxx} : dec_alu_input20_adrstage = 4'h4;  /* AND,A,B */
                    {8'h5c,2'bxx} : dec_alu_input20_adrstage = 4'h7;  /* AND,A,E */
                    {8'h5d,2'bxx} : dec_alu_input20_adrstage = 4'h6;  /* AND,A,D */
                    {8'h5e,2'bxx} : dec_alu_input20_adrstage = 4'h9;  /* AND,A,L */
                    {8'h5f,2'bxx} : dec_alu_input20_adrstage = 4'h8;  /* AND,A,H */
                    {8'h50,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* AND,X,A */
                    {8'h51,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* AND,A,A */
                    {8'h52,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* AND,C,A */
                    {8'h53,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* AND,B,A */
                    {8'h54,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* AND,E,A */
                    {8'h55,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* AND,D,A */
                    {8'h56,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* AND,L,A */
                    {8'h57,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* AND,H,A */
                    {8'hd0,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* AND,A,[HL+B] */
                    {8'hd2,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* AND,A,[HL+C] */
                    {8'h68,2'bxx} : dec_alu_input20_adrstage = 4'h3;  /* OR,A,X */
                    {8'h6a,2'bxx} : dec_alu_input20_adrstage = 4'h5;  /* OR,A,C */
                    {8'h6b,2'bxx} : dec_alu_input20_adrstage = 4'h4;  /* OR,A,B */
                    {8'h6c,2'bxx} : dec_alu_input20_adrstage = 4'h7;  /* OR,A,E */
                    {8'h6d,2'bxx} : dec_alu_input20_adrstage = 4'h6;  /* OR,A,D */
                    {8'h6e,2'bxx} : dec_alu_input20_adrstage = 4'h9;  /* OR,A,L */
                    {8'h6f,2'bxx} : dec_alu_input20_adrstage = 4'h8;  /* OR,A,H */
                    {8'h60,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* OR,X,A */
                    {8'h61,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* OR,A,A */
                    {8'h62,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* OR,C,A */
                    {8'h63,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* OR,B,A */
                    {8'h64,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* OR,E,A */
                    {8'h65,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* OR,D,A */
                    {8'h66,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* OR,L,A */
                    {8'h67,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* OR,H,A */
                    {8'he0,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* OR,A,[HL+B] */
                    {8'he2,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* OR,A,[HL+C] */
                    {8'h78,2'bxx} : dec_alu_input20_adrstage = 4'h3;  /* XOR,A,X */
                    {8'h7a,2'bxx} : dec_alu_input20_adrstage = 4'h5;  /* XOR,A,C */
                    {8'h7b,2'bxx} : dec_alu_input20_adrstage = 4'h4;  /* XOR,A,B */
                    {8'h7c,2'bxx} : dec_alu_input20_adrstage = 4'h7;  /* XOR,A,E */
                    {8'h7d,2'bxx} : dec_alu_input20_adrstage = 4'h6;  /* XOR,A,D */
                    {8'h7e,2'bxx} : dec_alu_input20_adrstage = 4'h9;  /* XOR,A,L */
                    {8'h7f,2'bxx} : dec_alu_input20_adrstage = 4'h8;  /* XOR,A,H */
                    {8'h70,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* XOR,X,A */
                    {8'h71,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* XOR,A,A */
                    {8'h72,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* XOR,C,A */
                    {8'h73,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* XOR,B,A */
                    {8'h74,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* XOR,E,A */
                    {8'h75,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* XOR,D,A */
                    {8'h76,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* XOR,L,A */
                    {8'h77,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* XOR,H,A */
                    {8'hf0,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* XOR,A,[HL+B] */
                    {8'hf2,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* XOR,A,[HL+C] */
                    {8'h48,2'bxx} : dec_alu_input20_adrstage = 4'h3;  /* CMP,A,X */
                    {8'h4a,2'bxx} : dec_alu_input20_adrstage = 4'h5;  /* CMP,A,C */
                    {8'h4b,2'bxx} : dec_alu_input20_adrstage = 4'h4;  /* CMP,A,B */
                    {8'h4c,2'bxx} : dec_alu_input20_adrstage = 4'h7;  /* CMP,A,E */
                    {8'h4d,2'bxx} : dec_alu_input20_adrstage = 4'h6;  /* CMP,A,D */
                    {8'h4e,2'bxx} : dec_alu_input20_adrstage = 4'h9;  /* CMP,A,L */
                    {8'h4f,2'bxx} : dec_alu_input20_adrstage = 4'h8;  /* CMP,A,H */
                    {8'h40,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* CMP,X,A */
                    {8'h41,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* CMP,A,A */
                    {8'h42,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* CMP,C,A */
                    {8'h43,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* CMP,B,A */
                    {8'h44,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* CMP,E,A */
                    {8'h45,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* CMP,D,A */
                    {8'h46,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* CMP,L,A */
                    {8'h47,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* CMP,H,A */
                    {8'hc0,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* CMP,A,[HL+B] */
                    {8'hc2,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* CMP,A,[HL+C] */
                    {8'hde,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* CMPS,X,[HL+byte] */
                    {8'h09,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* ADDW,AX,[HL+byte] */
                    {8'h29,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* SUBW,AX,[HL+byte] */
                    {8'h49,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* CMPW,AX,[HL+byte] */
                    {8'h59,2'bx0} : dec_alu_input20_adrstage = 4'h1;  /* INC,,[HL+byte] */
                    {8'h69,2'bx0} : dec_alu_input20_adrstage = 4'h1;  /* DEC,,[HL+byte] */
                    {8'h79,2'bx0} : dec_alu_input20_adrstage = 4'h1;  /* INCW,,[HL+byte] */
                    {8'h89,2'bx0} : dec_alu_input20_adrstage = 4'h1;  /* DECW,,[HL+byte] */
                    {8'hec,2'b00} : dec_alu_input20_adrstage = 4'hc;  /* RETB,, */
                    {8'hec,2'b01} : dec_alu_input20_adrstage = 4'hc;  /* RETB,, */
                    {8'hfc,2'b00} : dec_alu_input20_adrstage = 4'hc;  /* RETI,, */
                    {8'hfc,2'b01} : dec_alu_input20_adrstage = 4'hc;  /* RETI,, */
                    {8'hcd,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* POP,,PSW */
                    {8'hcf,2'bxx} : dec_alu_input20_adrstage = 4'ha;  /* SEL,,RB0 */
                    {8'hdf,2'bxx} : dec_alu_input20_adrstage = 4'ha;  /* SEL,,RB1 */
                    {8'hef,2'bxx} : dec_alu_input20_adrstage = 4'ha;  /* SEL,,RB2 */
                    {8'hff,2'bxx} : dec_alu_input20_adrstage = 4'ha;  /* SEL,,RB3 */
                    {8'h19,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* ADDC,A,A */
                    {8'h39,2'bxx} : dec_alu_input20_adrstage = 4'h2;  /* SUBC,A,A */
                    {8'hd1,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* AND,A,[HL+B] */
                    {8'he1,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* OR,A,[HL+B] */
                    {8'hf1,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* XOR,A,[HL+B] */
                    {8'h83,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* ADD,A,[HL+C] */
                    {8'h93,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* ADDC,A,[HL+C] */
                    {8'ha3,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* SUB,A,[HL+C] */
                    {8'hb3,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* SUBC,A,[HL+C] */
                    default : dec_alu_input20_adrstage = 4'h0;
                endcase
            end else if(ID_stage0 == 8'h71) begin
                    dec_alu_input20_adrstage = 4'h0;
            end else if(ID_stage0 == 8'h31) begin
                    dec_alu_input20_adrstage = 4'h0;
            end else begin
                casex ({ID_stage0,stage_adr})  
                    {8'h0c,2'bxx} : dec_alu_input20_adrstage = 4'ha;  /* ADD,A,#byte */
                    {8'h0a,2'bx0} : dec_alu_input20_adrstage = 4'ha;  /* ADD,saddr,#byte */
                    {8'h0b,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* ADD,A,saddr */
                    {8'h0f,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* ADD,A,!addr16 */
                    {8'h0d,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* ADD,A,[HL] */
                    {8'h0e,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* ADD,A,[HL+byte] */
                    {8'h1c,2'bxx} : dec_alu_input20_adrstage = 4'ha;  /* ADDC,A,#byte */
                    {8'h1a,2'bx0} : dec_alu_input20_adrstage = 4'ha;  /* ADDC,saddr,#byte */
                    {8'h1b,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* ADDC,A,saddr */
                    {8'h1f,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* ADDC,A,!addr16 */
                    {8'h1d,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* ADDC,A,[HL] */
                    {8'h1e,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* ADDC,A,[HL+byte] */
                    {8'h2c,2'bxx} : dec_alu_input20_adrstage = 4'ha;  /* SUB,A,#byte */
                    {8'h2a,2'bx0} : dec_alu_input20_adrstage = 4'ha;  /* SUB,saddr,#byte */
                    {8'h2b,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* SUB,A,saddr */
                    {8'h2f,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* SUB,A,!addr16 */
                    {8'h2d,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* SUB,A,[HL] */
                    {8'h2e,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* SUB,A,[HL+byte] */
                    {8'h3c,2'bxx} : dec_alu_input20_adrstage = 4'ha;  /* SUBC,A,#byte */
                    {8'h3a,2'bx0} : dec_alu_input20_adrstage = 4'ha;  /* SUBC,saddr,#byte */
                    {8'h3b,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* SUBC,A,saddr */
                    {8'h3f,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* SUBC,A,!addr16 */
                    {8'h3d,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* SUBC,A,[HL] */
                    {8'h3e,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* SUBC,A,[HL+byte] */
                    {8'h5c,2'bxx} : dec_alu_input20_adrstage = 4'ha;  /* AND,A,#byte */
                    {8'h5a,2'bx0} : dec_alu_input20_adrstage = 4'ha;  /* AND,saddr,#byte */
                    {8'h5b,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* AND,A,saddr */
                    {8'h5f,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* AND,A,!addr16 */
                    {8'h5d,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* AND,A,[HL] */
                    {8'h5e,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* AND,A,[HL+byte] */
                    {8'h6c,2'bxx} : dec_alu_input20_adrstage = 4'ha;  /* OR,A,#byte */
                    {8'h6a,2'bx0} : dec_alu_input20_adrstage = 4'ha;  /* OR,saddr,#byte */
                    {8'h6b,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* OR,A,saddr */
                    {8'h6f,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* OR,A,!addr16 */
                    {8'h6d,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* OR,A,[HL] */
                    {8'h6e,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* OR,A,[HL+byte] */
                    {8'h7c,2'bxx} : dec_alu_input20_adrstage = 4'ha;  /* XOR,A,#byte */
                    {8'h7a,2'bx0} : dec_alu_input20_adrstage = 4'ha;  /* XOR,saddr,#byte */
                    {8'h7b,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* XOR,A,saddr */
                    {8'h7f,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* XOR,A,!addr16 */
                    {8'h7d,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* XOR,A,[HL] */
                    {8'h7e,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* XOR,A,[HL+byte] */
                    {8'h4c,2'bxx} : dec_alu_input20_adrstage = 4'ha;  /* CMP,A,#byte */
                    {8'h4a,2'bxx} : dec_alu_input20_adrstage = 4'ha;  /* CMP,saddr,#byte */
                    {8'h40,2'bxx} : dec_alu_input20_adrstage = 4'ha;  /* CMP,!addr16,#byte */
                    {8'h4b,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* CMP,A,saddr */
                    {8'h4f,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* CMP,A,!addr16 */
                    {8'h4d,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* CMP,A,[HL] */
                    {8'h4e,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* CMP,A,[HL+byte] */
                    {8'h04,2'bxx} : dec_alu_input20_adrstage = 4'ha;  /* ADDW,AX,#word */
                    {8'h01,2'bxx} : dec_alu_input20_adrstage = 4'h3;  /* ADDW,AX,AX */
                    {8'h03,2'bxx} : dec_alu_input20_adrstage = 4'h5;  /* ADDW,AX,BC */
                    {8'h05,2'bxx} : dec_alu_input20_adrstage = 4'h7;  /* ADDW,AX,DE */
                    {8'h07,2'bxx} : dec_alu_input20_adrstage = 4'h9;  /* ADDW,AX,HL */
                    {8'h06,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* ADDW,AX,saddrp */
                    {8'h02,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* ADDW,AX,!addr16 */
                    {8'h24,2'bxx} : dec_alu_input20_adrstage = 4'ha;  /* SUBW,AX,#word */
                    {8'h21,2'bxx} : dec_alu_input20_adrstage = 4'h3;  /* SUBW,AX,AX */
                    {8'h23,2'bxx} : dec_alu_input20_adrstage = 4'h5;  /* SUBW,AX,BC */
                    {8'h25,2'bxx} : dec_alu_input20_adrstage = 4'h7;  /* SUBW,AX,DE */
                    {8'h27,2'bxx} : dec_alu_input20_adrstage = 4'h9;  /* SUBW,AX,HL */
                    {8'h26,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* SUBW,AX,saddrp */
                    {8'h22,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* SUBW,AX,!addr16 */
                    {8'h44,2'bxx} : dec_alu_input20_adrstage = 4'ha;  /* CMPW,AX,#word */
                    {8'h43,2'bxx} : dec_alu_input20_adrstage = 4'h5;  /* CMPW,AX,BC */
                    {8'h45,2'bxx} : dec_alu_input20_adrstage = 4'h7;  /* CMPW,AX,DE */
                    {8'h47,2'bxx} : dec_alu_input20_adrstage = 4'h9;  /* CMPW,AX,HL */
                    {8'h46,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* CMPW,AX,saddrp */
                    {8'h42,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* CMPW,AX,!addr16 */
                    {8'h80,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* INC,,X */
                    {8'h81,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* INC,,A */
                    {8'h82,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* INC,,C */
                    {8'h83,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* INC,,B */
                    {8'h84,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* INC,,E */
                    {8'h85,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* INC,,D */
                    {8'h86,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* INC,,L */
                    {8'h87,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* INC,,H */
                    {8'ha4,2'bx0} : dec_alu_input20_adrstage = 4'h1;  /* INC,,saddr */
                    {8'ha0,2'bx0} : dec_alu_input20_adrstage = 4'h1;  /* INC,,!addr16 */
                    {8'h90,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* DEC,,X */
                    {8'h91,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* DEC,,A */
                    {8'h92,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* DEC,,C */
                    {8'h93,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* DEC,,B */
                    {8'h94,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* DEC,,E */
                    {8'h95,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* DEC,,D */
                    {8'h96,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* DEC,,L */
                    {8'h97,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* DEC,,H */
                    {8'hb4,2'bx0} : dec_alu_input20_adrstage = 4'h1;  /* DEC,,saddr */
                    {8'hb0,2'bx0} : dec_alu_input20_adrstage = 4'h1;  /* DEC,,!addr16 */
                    {8'ha1,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* INCW,,AX */
                    {8'ha3,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* INCW,,BC */
                    {8'ha5,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* INCW,,DE */
                    {8'ha7,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* INCW,,HL */
                    {8'ha6,2'bx0} : dec_alu_input20_adrstage = 4'h1;  /* INCW,,saddrp */
                    {8'ha2,2'bx0} : dec_alu_input20_adrstage = 4'h1;  /* INCW,,!addr16 */
                    {8'hb1,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* DECW,,AX */
                    {8'hb3,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* DECW,,BC */
                    {8'hb5,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* DECW,,DE */
                    {8'hb7,2'bxx} : dec_alu_input20_adrstage = 4'h1;  /* DECW,,HL */
                    {8'hb6,2'bx0} : dec_alu_input20_adrstage = 4'h1;  /* DECW,,saddrp */
                    {8'hb2,2'bx0} : dec_alu_input20_adrstage = 4'h1;  /* DECW,,!addr16 */
                    {8'hd7,2'b00} : dec_alu_input20_adrstage = 4'hc;  /* RET,, */
                    {8'hd7,2'b01} : dec_alu_input20_adrstage = 4'hc;  /* RET,, */
                    {8'hc0,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* POP,,AX */
                    {8'hc2,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* POP,,BC */
                    {8'hc4,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* POP,,DE */
                    {8'hc6,2'bxx} : dec_alu_input20_adrstage = 4'hc;  /* POP,,HL */
                    {8'h10,2'bxx} : dec_alu_input20_adrstage = 4'hb;  /* ADDW,SP,#byte */
                    {8'h20,2'bxx} : dec_alu_input20_adrstage = 4'hb;  /* SUBW,SP,#byte */
                    default : dec_alu_input20_adrstage = 4'h0;
                endcase
            end
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_alu_input20 <= 4'h0;
        else if(cpuen) dec_alu_input20 <= dec_alu_input20_adrstage;
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*����INC,INCW,ADD,ADDC�Υ��ꥢ�������黻�򣲥���å��ܤ��飱����å��ܤ��ѹ�	*/
/*------------------------------------------------------------------------------*/

    output dec_alu_add;
    reg    dec_alu_add, dec_alu_add_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_alu_add_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h0c,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,A,#byte */
                {8'h0a,8'hxx,2'bx0} : dec_alu_add_adrstage = 1'b1;  /* ADD,saddr,#byte */
                {8'h61,8'h08,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,A,X */
                {8'h61,8'h0a,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,A,C */
                {8'h61,8'h0b,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,A,B */
                {8'h61,8'h0c,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,A,E */
                {8'h61,8'h0d,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,A,D */
                {8'h61,8'h0e,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,A,L */
                {8'h61,8'h0f,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,A,H */
                {8'h61,8'h00,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,X,A */
                {8'h61,8'h01,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,A,A */
                {8'h61,8'h02,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,C,A */
                {8'h61,8'h03,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,B,A */
                {8'h61,8'h04,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,E,A */
                {8'h61,8'h05,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,D,A */
                {8'h61,8'h06,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,L,A */
                {8'h61,8'h07,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,H,A */
                {8'h0b,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,A,saddr */
                {8'h0f,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,A,!addr16 */
                {8'h0d,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,A,[HL] */
                {8'h0e,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,A,[HL+byte] */
                {8'h61,8'h80,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,A,[HL+B] */
                {8'h61,8'h82,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,A,[HL+C] */
                {8'h1c,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,A,#byte */
                {8'h1a,8'hxx,2'bx0} : dec_alu_add_adrstage = 1'b1;  /* ADDC,saddr,#byte */
                {8'h61,8'h18,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,A,X */
                {8'h61,8'h1a,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,A,C */
                {8'h61,8'h1b,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,A,B */
                {8'h61,8'h1c,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,A,E */
                {8'h61,8'h1d,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,A,D */
                {8'h61,8'h1e,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,A,L */
                {8'h61,8'h1f,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,A,H */
                {8'h61,8'h10,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,X,A */
                {8'h61,8'h11,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,A,A */
                {8'h61,8'h12,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,C,A */
                {8'h61,8'h13,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,B,A */
                {8'h61,8'h14,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,E,A */
                {8'h61,8'h15,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,D,A */
                {8'h61,8'h16,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,L,A */
                {8'h61,8'h17,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,H,A */
                {8'h1b,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,A,saddr */
                {8'h1f,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,A,!addr16 */
                {8'h1d,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,A,[HL] */
                {8'h1e,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,A,[HL+byte] */
                {8'h61,8'h90,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,A,[HL+B] */
                {8'h61,8'h92,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,A,[HL+C] */
                {8'h04,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDW,AX,#word */
                {8'h01,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDW,AX,AX */
                {8'h03,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDW,AX,BC */
                {8'h05,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDW,AX,DE */
                {8'h07,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDW,AX,HL */
                {8'h06,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDW,AX,saddrp */
                {8'h02,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDW,AX,!addr16 */
                {8'h61,8'h09,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDW,AX,[HL+byte] */
                {8'h80,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* INC,,X */
                {8'h81,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* INC,,A */
                {8'h82,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* INC,,C */
                {8'h83,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* INC,,B */
                {8'h84,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* INC,,E */
                {8'h85,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* INC,,D */
                {8'h86,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* INC,,L */
                {8'h87,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* INC,,H */
                {8'ha4,8'hxx,2'bx0} : dec_alu_add_adrstage = 1'b1;  /* INC,,saddr */
                {8'ha0,8'hxx,2'bx0} : dec_alu_add_adrstage = 1'b1;  /* INC,,!addr16 */
                {8'h61,8'h59,2'bx0} : dec_alu_add_adrstage = 1'b1;  /* INC,,[HL+byte] */
                {8'ha1,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* INCW,,AX */
                {8'ha3,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* INCW,,BC */
                {8'ha5,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* INCW,,DE */
                {8'ha7,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* INCW,,HL */
                {8'ha6,8'hxx,2'bx0} : dec_alu_add_adrstage = 1'b1;  /* INCW,,saddrp */
                {8'ha2,8'hxx,2'bx0} : dec_alu_add_adrstage = 1'b1;  /* INCW,,!addr16 */
                {8'h61,8'h79,2'bx0} : dec_alu_add_adrstage = 1'b1;  /* INCW,,[HL+byte] */
                {8'h10,8'hxx,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDW,SP,#byte */
                {8'h61,8'h19,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,A,A */
                {8'h61,8'h83,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADD,A,[HL+C] */
                {8'h61,8'h93,2'bxx} : dec_alu_add_adrstage = 1'b1;  /* ADDC,A,[HL+C] */
                default : dec_alu_add_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_alu_add <= 1'b0;
        else if(cpuen) dec_alu_add <= dec_alu_add_adrstage;
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*����DEC,DECW,SUB,SUBC�Υ��ꥢ�������黻�򣲥���å��ܤ��飱����å��ܤ��ѹ�	*/
/*------------------------------------------------------------------------------*/

    output dec_alu_sub;
    reg    dec_alu_sub, dec_alu_sub_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_alu_sub_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h2c,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,A,#byte */
                {8'h2a,8'hxx,2'bx0} : dec_alu_sub_adrstage = 1'b1;  /* SUB,saddr,#byte */
                {8'h61,8'h28,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,A,X */
                {8'h61,8'h2a,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,A,C */
                {8'h61,8'h2b,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,A,B */
                {8'h61,8'h2c,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,A,E */
                {8'h61,8'h2d,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,A,D */
                {8'h61,8'h2e,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,A,L */
                {8'h61,8'h2f,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,A,H */
                {8'h61,8'h20,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,X,A */
                {8'h61,8'h21,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,A,A */
                {8'h61,8'h22,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,C,A */
                {8'h61,8'h23,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,B,A */
                {8'h61,8'h24,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,E,A */
                {8'h61,8'h25,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,D,A */
                {8'h61,8'h26,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,L,A */
                {8'h61,8'h27,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,H,A */
                {8'h2b,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,A,saddr */
                {8'h2f,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,A,!addr16 */
                {8'h2d,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,A,[HL] */
                {8'h2e,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,A,[HL+byte] */
                {8'h61,8'ha0,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,A,[HL+B] */
                {8'h61,8'ha2,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,A,[HL+C] */
                {8'h3c,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,A,#byte */
                {8'h3a,8'hxx,2'bx0} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,saddr,#byte */
                {8'h61,8'h38,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,A,X */
                {8'h61,8'h3a,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,A,C */
                {8'h61,8'h3b,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,A,B */
                {8'h61,8'h3c,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,A,E */
                {8'h61,8'h3d,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,A,D */
                {8'h61,8'h3e,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,A,L */
                {8'h61,8'h3f,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,A,H */
                {8'h61,8'h30,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,X,A */
                {8'h61,8'h31,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,A,A */
                {8'h61,8'h32,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,C,A */
                {8'h61,8'h33,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,B,A */
                {8'h61,8'h34,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,E,A */
                {8'h61,8'h35,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,D,A */
                {8'h61,8'h36,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,L,A */
                {8'h61,8'h37,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,H,A */
                {8'h3b,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,A,saddr */
                {8'h3f,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,A,!addr16 */
                {8'h3d,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,A,[HL] */
                {8'h3e,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,A,[HL+byte] */
                {8'h61,8'hb0,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,A,[HL+B] */
                {8'h61,8'hb2,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,A,[HL+C] */
                {8'h4c,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,A,#byte */
                {8'h4a,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,saddr,#byte */
                {8'h40,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,!addr16,#byte */
                {8'h61,8'h48,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,A,X */
                {8'h61,8'h4a,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,A,C */
                {8'h61,8'h4b,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,A,B */
                {8'h61,8'h4c,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,A,E */
                {8'h61,8'h4d,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,A,D */
                {8'h61,8'h4e,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,A,L */
                {8'h61,8'h4f,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,A,H */
                {8'h61,8'h40,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,X,A */
                {8'h61,8'h41,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,A,A */
                {8'h61,8'h42,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,C,A */
                {8'h61,8'h43,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,B,A */
                {8'h61,8'h44,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,E,A */
                {8'h61,8'h45,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,D,A */
                {8'h61,8'h46,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,L,A */
                {8'h61,8'h47,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,H,A */
                {8'h4b,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,A,saddr */
                {8'h4f,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,A,!addr16 */
                {8'h4d,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,A,[HL] */
                {8'h4e,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,A,[HL+byte] */
                {8'h61,8'hc0,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,A,[HL+B] */
                {8'h61,8'hc2,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP,A,[HL+C] */
                {8'h61,8'hde,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMPS,X,[HL+byte] */
                {8'hd1,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP0,,A */
                {8'hd0,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP0,,X */
                {8'hd3,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP0,,B */
                {8'hd2,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP0,,C */
                {8'hd4,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP0,,saddr */
                {8'hd5,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMP0,,!addr16 */
                {8'h24,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBW,AX,#word */
                {8'h21,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBW,AX,AX */
                {8'h23,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBW,AX,BC */
                {8'h25,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBW,AX,DE */
                {8'h27,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBW,AX,HL */
                {8'h26,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBW,AX,saddrp */
                {8'h22,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBW,AX,!addr16 */
                {8'h61,8'h29,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBW,AX,[HL+byte] */
                {8'h44,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMPW,AX,#word */
                {8'h43,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMPW,AX,BC */
                {8'h45,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMPW,AX,DE */
                {8'h47,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMPW,AX,HL */
                {8'h46,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMPW,AX,saddrp */
                {8'h42,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMPW,AX,!addr16 */
                {8'h61,8'h49,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* CMPW,AX,[HL+byte] */
                {8'h90,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* DEC,,X */
                {8'h91,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* DEC,,A */
                {8'h92,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* DEC,,C */
                {8'h93,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* DEC,,B */
                {8'h94,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* DEC,,E */
                {8'h95,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* DEC,,D */
                {8'h96,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* DEC,,L */
                {8'h97,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* DEC,,H */
                {8'hb4,8'hxx,2'bx0} : dec_alu_sub_adrstage = 1'b1;  /* DEC,,saddr */
                {8'hb0,8'hxx,2'bx0} : dec_alu_sub_adrstage = 1'b1;  /* DEC,,!addr16 */
                {8'h61,8'h69,2'bx0} : dec_alu_sub_adrstage = 1'b1;  /* DEC,,[HL+byte] */
                {8'hb1,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* DECW,,AX */
                {8'hb3,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* DECW,,BC */
                {8'hb5,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* DECW,,DE */
                {8'hb7,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* DECW,,HL */
                {8'hb6,8'hxx,2'bx0} : dec_alu_sub_adrstage = 1'b1;  /* DECW,,saddrp */
                {8'hb2,8'hxx,2'bx0} : dec_alu_sub_adrstage = 1'b1;  /* DECW,,!addr16 */
                {8'h61,8'h89,2'bx0} : dec_alu_sub_adrstage = 1'b1;  /* DECW,,[HL+byte] */
                {8'h20,8'hxx,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBW,SP,#byte */
                {8'h61,8'h39,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,A,A */
                {8'h61,8'ha3,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUB,A,[HL+C] */
                {8'h61,8'hb3,2'bxx} : dec_alu_sub_adrstage = 1'b1;  /* SUBC,A,[HL+C] */
                default : dec_alu_sub_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_alu_sub <= 1'b0;
        else if(cpuen) dec_alu_sub <= dec_alu_sub_adrstage;
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*����AND�Υ��ꥢ�������黻�򣲥���å��ܤ��飱����å��ܤ��ѹ�		*/
/*����AND1,CLR1,BTCLR�����̺����dec_alu_andbit�ذ�ư				*/
/*------------------------------------------------------------------------------*/

    output dec_alu_and;
    reg    dec_alu_and, dec_alu_and_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_alu_and_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h5c,8'hxx,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,A,#byte */
                {8'h5a,8'hxx,2'bx0} : dec_alu_and_adrstage = 1'b1;  /* AND,saddr,#byte */
                {8'h61,8'h58,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,A,X */
                {8'h61,8'h5a,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,A,C */
                {8'h61,8'h5b,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,A,B */
                {8'h61,8'h5c,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,A,E */
                {8'h61,8'h5d,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,A,D */
                {8'h61,8'h5e,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,A,L */
                {8'h61,8'h5f,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,A,H */
                {8'h61,8'h50,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,X,A */
                {8'h61,8'h51,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,A,A */
                {8'h61,8'h52,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,C,A */
                {8'h61,8'h53,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,B,A */
                {8'h61,8'h54,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,E,A */
                {8'h61,8'h55,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,D,A */
                {8'h61,8'h56,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,L,A */
                {8'h61,8'h57,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,H,A */
                {8'h5b,8'hxx,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,A,saddr */
                {8'h5f,8'hxx,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,A,!addr16 */
                {8'h5d,8'hxx,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,A,[HL] */
                {8'h5e,8'hxx,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,A,[HL+byte] */
                {8'h61,8'hd0,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,A,[HL+B] */
                {8'h61,8'hd2,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,A,[HL+C] */
                {8'h61,8'hd1,2'bxx} : dec_alu_and_adrstage = 1'b1;  /* AND,A,[HL+B] */
                default : dec_alu_and_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_alu_and <= 1'b0;
        else if(cpuen) dec_alu_and <= dec_alu_and_adrstage;
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ӥå����̿��(AND1,CLR1,BTCLR)�����Ѳ�					*/
/*------------------------------------------------------------------------------*/

    output dec_alu_andbit;
    reg    dec_alu_andbit, dec_alu_andbit_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_alu_andbit_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h71,8'h05,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,saddr.0 */
                {8'h71,8'h15,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,saddr.1 */
                {8'h71,8'h25,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,saddr.2 */
                {8'h71,8'h35,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,saddr.3 */
                {8'h71,8'h45,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,saddr.4 */
                {8'h71,8'h55,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,saddr.5 */
                {8'h71,8'h65,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,saddr.6 */
                {8'h71,8'h75,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,saddr.7 */
                {8'h71,8'h0d,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,sfr.0 */
                {8'h71,8'h1d,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,sfr.1 */
                {8'h71,8'h2d,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,sfr.2 */
                {8'h71,8'h3d,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,sfr.3 */
                {8'h71,8'h4d,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,sfr.4 */
                {8'h71,8'h5d,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,sfr.5 */
                {8'h71,8'h6d,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,sfr.6 */
                {8'h71,8'h7d,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,sfr.7 */
                {8'h71,8'h8d,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,A.0 */
                {8'h71,8'h9d,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,A.1 */
                {8'h71,8'had,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,A.2 */
                {8'h71,8'hbd,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,A.3 */
                {8'h71,8'hcd,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,A.4 */
                {8'h71,8'hdd,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,A.5 */
                {8'h71,8'hed,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,A.6 */
                {8'h71,8'hfd,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,A.7 */
                {8'h71,8'h85,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,[HL].0 */
                {8'h71,8'h95,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,[HL].1 */
                {8'h71,8'ha5,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,[HL].2 */
                {8'h71,8'hb5,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,[HL].3 */
                {8'h71,8'hc5,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,[HL].4 */
                {8'h71,8'hd5,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,[HL].5 */
                {8'h71,8'he5,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,[HL].6 */
                {8'h71,8'hf5,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* AND1,CY,[HL].7 */
                {8'h71,8'h03,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,saddr.0 */
                {8'h71,8'h13,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,saddr.1 */
                {8'h71,8'h23,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,saddr.2 */
                {8'h71,8'h33,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,saddr.3 */
                {8'h71,8'h43,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,saddr.4 */
                {8'h71,8'h53,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,saddr.5 */
                {8'h71,8'h63,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,saddr.6 */
                {8'h71,8'h73,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,saddr.7 */
                {8'h71,8'h0b,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,sfr.0 */
                {8'h71,8'h1b,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,sfr.1 */
                {8'h71,8'h2b,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,sfr.2 */
                {8'h71,8'h3b,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,sfr.3 */
                {8'h71,8'h4b,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,sfr.4 */
                {8'h71,8'h5b,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,sfr.5 */
                {8'h71,8'h6b,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,sfr.6 */
                {8'h71,8'h7b,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,sfr.7 */
                {8'h71,8'h8b,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,A.0 */
                {8'h71,8'h9b,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,A.1 */
                {8'h71,8'hab,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,A.2 */
                {8'h71,8'hbb,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,A.3 */
                {8'h71,8'hcb,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,A.4 */
                {8'h71,8'hdb,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,A.5 */
                {8'h71,8'heb,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,A.6 */
                {8'h71,8'hfb,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,A.7 */
                {8'h71,8'h08,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,!addr16.0 */
                {8'h71,8'h18,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,!addr16.1 */
                {8'h71,8'h28,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,!addr16.2 */
                {8'h71,8'h38,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,!addr16.3 */
                {8'h71,8'h48,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,!addr16.4 */
                {8'h71,8'h58,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,!addr16.5 */
                {8'h71,8'h68,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,!addr16.6 */
                {8'h71,8'h78,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,!addr16.7 */
                {8'h71,8'h83,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,[HL].0 */
                {8'h71,8'h93,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,[HL].1 */
                {8'h71,8'ha3,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,[HL].2 */
                {8'h71,8'hb3,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,[HL].3 */
                {8'h71,8'hc3,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,[HL].4 */
                {8'h71,8'hd3,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,[HL].5 */
                {8'h71,8'he3,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,[HL].6 */
                {8'h71,8'hf3,2'bx0} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,[HL].7 */
                {8'h71,8'h88,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,CY */
                {8'h71,8'h98,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,CY */
                {8'h71,8'ha8,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,CY */
                {8'h71,8'hb8,2'bxx} : dec_alu_andbit_adrstage = 1'b1;  /* CLR1,,CY */
                {8'h31,8'h00,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,saddr.0,$addr8 */
                {8'h31,8'h10,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,saddr.1,$addr8 */
                {8'h31,8'h20,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,saddr.2,$addr8 */
                {8'h31,8'h30,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,saddr.3,$addr8 */
                {8'h31,8'h40,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,saddr.4,$addr8 */
                {8'h31,8'h50,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,saddr.5,$addr8 */
                {8'h31,8'h60,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,saddr.6,$addr8 */
                {8'h31,8'h70,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,saddr.7,$addr8 */
                {8'h31,8'h80,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,sfr.0,$addr8 */
                {8'h31,8'h90,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,sfr.1,$addr8 */
                {8'h31,8'ha0,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,sfr.2,$addr8 */
                {8'h31,8'hb0,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,sfr.3,$addr8 */
                {8'h31,8'hc0,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,sfr.4,$addr8 */
                {8'h31,8'hd0,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,sfr.5,$addr8 */
                {8'h31,8'he0,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,sfr.6,$addr8 */
                {8'h31,8'hf0,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,sfr.7,$addr8 */
                {8'h31,8'h01,2'b10} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,A.0,$addr8 */
                {8'h31,8'h11,2'b10} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,A.1,$addr8 */
                {8'h31,8'h21,2'b10} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,A.2,$addr8 */
                {8'h31,8'h31,2'b10} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,A.3,$addr8 */
                {8'h31,8'h41,2'b10} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,A.4,$addr8 */
                {8'h31,8'h51,2'b10} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,A.5,$addr8 */
                {8'h31,8'h61,2'b10} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,A.6,$addr8 */
                {8'h31,8'h71,2'b10} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,A.7,$addr8 */
                {8'h31,8'h81,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,[HL].0,$addr8 */
                {8'h31,8'h91,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,[HL].1,$addr8 */
                {8'h31,8'ha1,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,[HL].2,$addr8 */
                {8'h31,8'hb1,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,[HL].3,$addr8 */
                {8'h31,8'hc1,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,[HL].4,$addr8 */
                {8'h31,8'hd1,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,[HL].5,$addr8 */
                {8'h31,8'he1,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,[HL].6,$addr8 */
                {8'h31,8'hf1,2'b01} : dec_alu_andbit_adrstage = 1'b1;  /* BTCLR,[HL].7,$addr8 */
                default : dec_alu_andbit_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_alu_andbit <= 1'b0;
        else if(cpuen) dec_alu_andbit <= dec_alu_andbit_adrstage;
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*����OR�Υ��ꥢ�������黻�򣲥���å��ܤ��飱����å��ܤ��ѹ�		*/
/*����OR1,SET1�����̺����dec_alu_orbit�ذ�ư					*/
/*����ONEB,ONEW�����̺����dec_alu_transout�ذ�ư				*/
/*------------------------------------------------------------------------------*/

    output dec_alu_or;
    reg    dec_alu_or, dec_alu_or_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_alu_or_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h6c,8'hxx,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,A,#byte */
                {8'h6a,8'hxx,2'bx0} : dec_alu_or_adrstage = 1'b1;  /* OR,saddr,#byte */
                {8'h61,8'h68,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,A,X */
                {8'h61,8'h6a,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,A,C */
                {8'h61,8'h6b,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,A,B */
                {8'h61,8'h6c,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,A,E */
                {8'h61,8'h6d,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,A,D */
                {8'h61,8'h6e,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,A,L */
                {8'h61,8'h6f,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,A,H */
                {8'h61,8'h60,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,X,A */
                {8'h61,8'h61,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,A,A */
                {8'h61,8'h62,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,C,A */
                {8'h61,8'h63,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,B,A */
                {8'h61,8'h64,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,E,A */
                {8'h61,8'h65,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,D,A */
                {8'h61,8'h66,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,L,A */
                {8'h61,8'h67,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,H,A */
                {8'h6b,8'hxx,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,A,saddr */
                {8'h6f,8'hxx,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,A,!addr16 */
                {8'h6d,8'hxx,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,A,[HL] */
                {8'h6e,8'hxx,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,A,[HL+byte] */
                {8'h61,8'he0,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,A,[HL+B] */
                {8'h61,8'he2,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,A,[HL+C] */
                {8'h61,8'he1,2'bxx} : dec_alu_or_adrstage = 1'b1;  /* OR,A,[HL+B] */
                default : dec_alu_or_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_alu_or <= 1'b0;
        else if(cpuen) dec_alu_or <= dec_alu_or_adrstage;
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ӥå����̿��(OR1,SET1)�����Ѳ�						*/
/*------------------------------------------------------------------------------*/

    output dec_alu_orbit;
    reg    dec_alu_orbit, dec_alu_orbit_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_alu_orbit_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h71,8'h06,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,saddr.0 */
                {8'h71,8'h16,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,saddr.1 */
                {8'h71,8'h26,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,saddr.2 */
                {8'h71,8'h36,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,saddr.3 */
                {8'h71,8'h46,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,saddr.4 */
                {8'h71,8'h56,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,saddr.5 */
                {8'h71,8'h66,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,saddr.6 */
                {8'h71,8'h76,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,saddr.7 */
                {8'h71,8'h0e,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,sfr.0 */
                {8'h71,8'h1e,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,sfr.1 */
                {8'h71,8'h2e,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,sfr.2 */
                {8'h71,8'h3e,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,sfr.3 */
                {8'h71,8'h4e,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,sfr.4 */
                {8'h71,8'h5e,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,sfr.5 */
                {8'h71,8'h6e,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,sfr.6 */
                {8'h71,8'h7e,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,sfr.7 */
                {8'h71,8'h8e,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,A.0 */
                {8'h71,8'h9e,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,A.1 */
                {8'h71,8'hae,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,A.2 */
                {8'h71,8'hbe,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,A.3 */
                {8'h71,8'hce,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,A.4 */
                {8'h71,8'hde,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,A.5 */
                {8'h71,8'hee,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,A.6 */
                {8'h71,8'hfe,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,A.7 */
                {8'h71,8'h86,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,[HL].0 */
                {8'h71,8'h96,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,[HL].1 */
                {8'h71,8'ha6,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,[HL].2 */
                {8'h71,8'hb6,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,[HL].3 */
                {8'h71,8'hc6,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,[HL].4 */
                {8'h71,8'hd6,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,[HL].5 */
                {8'h71,8'he6,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,[HL].6 */
                {8'h71,8'hf6,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* OR1,CY,[HL].7 */
                {8'h71,8'h02,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,saddr.0 */
                {8'h71,8'h12,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,saddr.1 */
                {8'h71,8'h22,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,saddr.2 */
                {8'h71,8'h32,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,saddr.3 */
                {8'h71,8'h42,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,saddr.4 */
                {8'h71,8'h52,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,saddr.5 */
                {8'h71,8'h62,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,saddr.6 */
                {8'h71,8'h72,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,saddr.7 */
                {8'h71,8'h0a,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,sfr.0 */
                {8'h71,8'h1a,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,sfr.1 */
                {8'h71,8'h2a,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,sfr.2 */
                {8'h71,8'h3a,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,sfr.3 */
                {8'h71,8'h4a,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,sfr.4 */
                {8'h71,8'h5a,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,sfr.5 */
                {8'h71,8'h6a,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,sfr.6 */
                {8'h71,8'h7a,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,sfr.7 */
                {8'h71,8'h8a,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,A.0 */
                {8'h71,8'h9a,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,A.1 */
                {8'h71,8'haa,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,A.2 */
                {8'h71,8'hba,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,A.3 */
                {8'h71,8'hca,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,A.4 */
                {8'h71,8'hda,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,A.5 */
                {8'h71,8'hea,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,A.6 */
                {8'h71,8'hfa,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,A.7 */
                {8'h71,8'h00,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,!addr16.0 */
                {8'h71,8'h10,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,!addr16.1 */
                {8'h71,8'h20,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,!addr16.2 */
                {8'h71,8'h30,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,!addr16.3 */
                {8'h71,8'h40,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,!addr16.4 */
                {8'h71,8'h50,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,!addr16.5 */
                {8'h71,8'h60,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,!addr16.6 */
                {8'h71,8'h70,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,!addr16.7 */
                {8'h71,8'h82,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,[HL].0 */
                {8'h71,8'h92,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,[HL].1 */
                {8'h71,8'ha2,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,[HL].2 */
                {8'h71,8'hb2,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,[HL].3 */
                {8'h71,8'hc2,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,[HL].4 */
                {8'h71,8'hd2,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,[HL].5 */
                {8'h71,8'he2,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,[HL].6 */
                {8'h71,8'hf2,2'bx0} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,[HL].7 */
                {8'h71,8'h80,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,CY */
                {8'h71,8'h90,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,CY */
                {8'h71,8'ha0,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,CY */
                {8'h71,8'hb0,2'bxx} : dec_alu_orbit_adrstage = 1'b1;  /* SET1,,CY */
                default : dec_alu_orbit_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_alu_orbit <= 1'b0;
        else if(cpuen) dec_alu_orbit <= dec_alu_orbit_adrstage;
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*����XOR�Υ��ꥢ�������黻�򣲥���å��ܤ��飱����å��ܤ��ѹ�		*/
/*����XOR1,BF,NOT1�����̺����dec_alu_andbit�ذ�ư				*/
/*------------------------------------------------------------------------------*/

    output dec_alu_exor;
    reg    dec_alu_exor, dec_alu_exor_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_alu_exor_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h7c,8'hxx,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,A,#byte */
                {8'h7a,8'hxx,2'bx0} : dec_alu_exor_adrstage = 1'b1;  /* XOR,saddr,#byte */
                {8'h61,8'h78,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,A,X */
                {8'h61,8'h7a,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,A,C */
                {8'h61,8'h7b,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,A,B */
                {8'h61,8'h7c,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,A,E */
                {8'h61,8'h7d,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,A,D */
                {8'h61,8'h7e,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,A,L */
                {8'h61,8'h7f,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,A,H */
                {8'h61,8'h70,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,X,A */
                {8'h61,8'h71,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,A,A */
                {8'h61,8'h72,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,C,A */
                {8'h61,8'h73,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,B,A */
                {8'h61,8'h74,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,E,A */
                {8'h61,8'h75,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,D,A */
                {8'h61,8'h76,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,L,A */
                {8'h61,8'h77,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,H,A */
                {8'h7b,8'hxx,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,A,saddr */
                {8'h7f,8'hxx,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,A,!addr16 */
                {8'h7d,8'hxx,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,A,[HL] */
                {8'h7e,8'hxx,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,A,[HL+byte] */
                {8'h61,8'hf0,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,A,[HL+B] */
                {8'h61,8'hf2,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,A,[HL+C] */
                {8'h61,8'hf1,2'bxx} : dec_alu_exor_adrstage = 1'b1;  /* XOR,A,[HL+B] */
                default : dec_alu_exor_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_alu_exor <= 1'b0;
        else if(cpuen) dec_alu_exor <= dec_alu_exor_adrstage;
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ӥå����̿��(XOR1,BF,NOT1)�����Ѳ�					*/
/*------------------------------------------------------------------------------*/

    output dec_alu_exorbit;
    reg    dec_alu_exorbit, dec_alu_exorbit_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_alu_exorbit_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h71,8'h07,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,saddr.0 */
                {8'h71,8'h17,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,saddr.1 */
                {8'h71,8'h27,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,saddr.2 */
                {8'h71,8'h37,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,saddr.3 */
                {8'h71,8'h47,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,saddr.4 */
                {8'h71,8'h57,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,saddr.5 */
                {8'h71,8'h67,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,saddr.6 */
                {8'h71,8'h77,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,saddr.7 */
                {8'h71,8'h0f,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,sfr.0 */
                {8'h71,8'h1f,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,sfr.1 */
                {8'h71,8'h2f,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,sfr.2 */
                {8'h71,8'h3f,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,sfr.3 */
                {8'h71,8'h4f,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,sfr.4 */
                {8'h71,8'h5f,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,sfr.5 */
                {8'h71,8'h6f,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,sfr.6 */
                {8'h71,8'h7f,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,sfr.7 */
                {8'h71,8'h8f,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,A.0 */
                {8'h71,8'h9f,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,A.1 */
                {8'h71,8'haf,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,A.2 */
                {8'h71,8'hbf,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,A.3 */
                {8'h71,8'hcf,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,A.4 */
                {8'h71,8'hdf,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,A.5 */
                {8'h71,8'hef,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,A.6 */
                {8'h71,8'hff,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,A.7 */
                {8'h71,8'h87,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,[HL].0 */
                {8'h71,8'h97,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,[HL].1 */
                {8'h71,8'ha7,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,[HL].2 */
                {8'h71,8'hb7,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,[HL].3 */
                {8'h71,8'hc7,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,[HL].4 */
                {8'h71,8'hd7,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,[HL].5 */
                {8'h71,8'he7,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,[HL].6 */
                {8'h71,8'hf7,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* XOR1,CY,[HL].7 */
                {8'h71,8'hc0,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* NOT1,,CY */
                {8'h71,8'hd0,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* NOT1,,CY */
                {8'h71,8'he0,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* NOT1,,CY */
                {8'h71,8'hf0,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* NOT1,,CY */
                {8'h71,8'hc8,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* NOT1,,CY */
                {8'h71,8'hd8,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* NOT1,,CY */
                {8'h71,8'he8,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* NOT1,,CY */
                {8'h71,8'hf8,2'bxx} : dec_alu_exorbit_adrstage = 1'b1;  /* NOT1,,CY */
                {8'h31,8'h04,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,saddr.0,$addr8 */
                {8'h31,8'h14,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,saddr.1,$addr8 */
                {8'h31,8'h24,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,saddr.2,$addr8 */
                {8'h31,8'h34,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,saddr.3,$addr8 */
                {8'h31,8'h44,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,saddr.4,$addr8 */
                {8'h31,8'h54,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,saddr.5,$addr8 */
                {8'h31,8'h64,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,saddr.6,$addr8 */
                {8'h31,8'h74,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,saddr.7,$addr8 */
                {8'h31,8'h84,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,sfr.0,$addr8 */
                {8'h31,8'h94,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,sfr.1,$addr8 */
                {8'h31,8'ha4,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,sfr.2,$addr8 */
                {8'h31,8'hb4,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,sfr.3,$addr8 */
                {8'h31,8'hc4,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,sfr.4,$addr8 */
                {8'h31,8'hd4,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,sfr.5,$addr8 */
                {8'h31,8'he4,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,sfr.6,$addr8 */
                {8'h31,8'hf4,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,sfr.7,$addr8 */
                {8'h31,8'h05,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,A.0,$addr8 */
                {8'h31,8'h15,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,A.1,$addr8 */
                {8'h31,8'h25,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,A.2,$addr8 */
                {8'h31,8'h35,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,A.3,$addr8 */
                {8'h31,8'h45,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,A.4,$addr8 */
                {8'h31,8'h55,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,A.5,$addr8 */
                {8'h31,8'h65,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,A.6,$addr8 */
                {8'h31,8'h75,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,A.7,$addr8 */
                {8'h31,8'h85,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,[HL].0,$addr8 */
                {8'h31,8'h95,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,[HL].1,$addr8 */
                {8'h31,8'ha5,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,[HL].2,$addr8 */
                {8'h31,8'hb5,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,[HL].3,$addr8 */
                {8'h31,8'hc5,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,[HL].4,$addr8 */
                {8'h31,8'hd5,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,[HL].5,$addr8 */
                {8'h31,8'he5,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,[HL].6,$addr8 */
                {8'h31,8'hf5,2'b00} : dec_alu_exorbit_adrstage = 1'b1;  /* BF,[HL].7,$addr8 */
                default : dec_alu_exorbit_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_alu_exorbit <= 1'b0;
        else if(cpuen) dec_alu_exorbit <= dec_alu_exorbit_adrstage;
    end

    output dec_alu_ror;
    reg    dec_alu_ror, dec_alu_ror_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_alu_ror_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hdb,2'bxx} : dec_alu_ror_adrstage = 1'b1;  /* ROR,A,1 */
                {8'h61,8'hfb,2'bxx} : dec_alu_ror_adrstage = 1'b1;  /* RORC,A,1 */
                default : dec_alu_ror_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_alu_ror <= 1'b0;
        else if(cpuen) dec_alu_ror <= dec_alu_ror_adrstage;
    end
    output dec_alu_rol;
    reg    dec_alu_rol, dec_alu_rol_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_alu_rol_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'heb,2'bxx} : dec_alu_rol_adrstage = 1'b1;  /* ROL,A,1 */
                {8'h61,8'hdc,2'bxx} : dec_alu_rol_adrstage = 1'b1;  /* ROLC,A,1 */
                {8'h61,8'hee,2'bxx} : dec_alu_rol_adrstage = 1'b1;  /* ROLWC,AX,1 */
                {8'h61,8'hfe,2'bxx} : dec_alu_rol_adrstage = 1'b1;  /* ROLWC,BC,1 */
                default : dec_alu_rol_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_alu_rol <= 1'b0;
        else if(cpuen) dec_alu_rol <= dec_alu_rol_adrstage;
    end
    output dec_alu_shr;
    reg    dec_alu_shr, dec_alu_shr_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_alu_shr_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h31,8'h0a,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHR,A,0 */
                {8'h31,8'h1a,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHR,A,1 */
                {8'h31,8'h2a,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHR,A,2 */
                {8'h31,8'h3a,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHR,A,3 */
                {8'h31,8'h4a,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHR,A,4 */
                {8'h31,8'h5a,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHR,A,5 */
                {8'h31,8'h6a,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHR,A,6 */
                {8'h31,8'h7a,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHR,A,7 */
                {8'h31,8'h0e,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHRW,AX,0 */
                {8'h31,8'h1e,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHRW,AX,1 */
                {8'h31,8'h2e,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHRW,AX,2 */
                {8'h31,8'h3e,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHRW,AX,3 */
                {8'h31,8'h4e,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHRW,AX,4 */
                {8'h31,8'h5e,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHRW,AX,5 */
                {8'h31,8'h6e,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHRW,AX,6 */
                {8'h31,8'h7e,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHRW,AX,7 */
                {8'h31,8'h8e,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHRW,AX,8 */
                {8'h31,8'h9e,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHRW,AX,9 */
                {8'h31,8'hae,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHRW,AX,10 */
                {8'h31,8'hbe,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHRW,AX,11 */
                {8'h31,8'hce,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHRW,AX,12 */
                {8'h31,8'hde,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHRW,AX,13 */
                {8'h31,8'hee,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHRW,AX,14 */
                {8'h31,8'hfe,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHRW,AX,15 */
                {8'h31,8'h8a,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHR,A,0 */
                {8'h31,8'h9a,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHR,A,1 */
                {8'h31,8'haa,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHR,A,2 */
                {8'h31,8'hba,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHR,A,3 */
                {8'h31,8'hca,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHR,A,4 */
                {8'h31,8'hda,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHR,A,5 */
                {8'h31,8'hea,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHR,A,6 */
                {8'h31,8'hfa,2'bxx} : dec_alu_shr_adrstage = 1'b1;  /* SHR,A,7 */
                default : dec_alu_shr_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_alu_shr <= 1'b0;
        else if(cpuen) dec_alu_shr <= dec_alu_shr_adrstage;
    end
    output dec_alu_shl;
    reg    dec_alu_shl, dec_alu_shl_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_alu_shl_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h31,8'h09,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,A,0 */
                {8'h31,8'h19,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,A,1 */
                {8'h31,8'h29,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,A,2 */
                {8'h31,8'h39,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,A,3 */
                {8'h31,8'h49,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,A,4 */
                {8'h31,8'h59,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,A,5 */
                {8'h31,8'h69,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,A,6 */
                {8'h31,8'h79,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,A,7 */
                {8'h31,8'h08,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,B,0 */
                {8'h31,8'h18,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,B,1 */
                {8'h31,8'h28,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,B,2 */
                {8'h31,8'h38,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,B,3 */
                {8'h31,8'h48,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,B,4 */
                {8'h31,8'h58,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,B,5 */
                {8'h31,8'h68,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,B,6 */
                {8'h31,8'h78,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,B,7 */
                {8'h31,8'h07,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,C,0 */
                {8'h31,8'h17,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,C,1 */
                {8'h31,8'h27,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,C,2 */
                {8'h31,8'h37,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,C,3 */
                {8'h31,8'h47,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,C,4 */
                {8'h31,8'h57,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,C,5 */
                {8'h31,8'h67,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,C,6 */
                {8'h31,8'h77,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,C,7 */
                {8'h31,8'h0d,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,AX,0 */
                {8'h31,8'h1d,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,AX,1 */
                {8'h31,8'h2d,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,AX,2 */
                {8'h31,8'h3d,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,AX,3 */
                {8'h31,8'h4d,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,AX,4 */
                {8'h31,8'h5d,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,AX,5 */
                {8'h31,8'h6d,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,AX,6 */
                {8'h31,8'h7d,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,AX,7 */
                {8'h31,8'h8d,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,AX,8 */
                {8'h31,8'h9d,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,AX,9 */
                {8'h31,8'had,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,AX,10 */
                {8'h31,8'hbd,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,AX,11 */
                {8'h31,8'hcd,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,AX,12 */
                {8'h31,8'hdd,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,AX,13 */
                {8'h31,8'hed,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,AX,14 */
                {8'h31,8'hfd,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,AX,15 */
                {8'h31,8'h0c,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,BC,0 */
                {8'h31,8'h1c,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,BC,1 */
                {8'h31,8'h2c,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,BC,2 */
                {8'h31,8'h3c,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,BC,3 */
                {8'h31,8'h4c,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,BC,4 */
                {8'h31,8'h5c,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,BC,5 */
                {8'h31,8'h6c,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,BC,6 */
                {8'h31,8'h7c,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,BC,7 */
                {8'h31,8'h8c,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,BC,8 */
                {8'h31,8'h9c,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,BC,9 */
                {8'h31,8'hac,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,BC,10 */
                {8'h31,8'hbc,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,BC,11 */
                {8'h31,8'hcc,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,BC,12 */
                {8'h31,8'hdc,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,BC,13 */
                {8'h31,8'hec,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,BC,14 */
                {8'h31,8'hfc,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHLW,BC,15 */
                {8'h31,8'h89,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,A,0 */
                {8'h31,8'h99,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,A,1 */
                {8'h31,8'ha9,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,A,2 */
                {8'h31,8'hb9,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,A,3 */
                {8'h31,8'hc9,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,A,4 */
                {8'h31,8'hd9,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,A,5 */
                {8'h31,8'he9,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,A,6 */
                {8'h31,8'hf9,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,A,7 */
                {8'h31,8'h88,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,B,0 */
                {8'h31,8'h98,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,B,1 */
                {8'h31,8'ha8,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,B,2 */
                {8'h31,8'hb8,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,B,3 */
                {8'h31,8'hc8,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,B,4 */
                {8'h31,8'hd8,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,B,5 */
                {8'h31,8'he8,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,B,6 */
                {8'h31,8'hf8,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,B,7 */
                {8'h31,8'h87,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,C,0 */
                {8'h31,8'h97,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,C,1 */
                {8'h31,8'ha7,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,C,2 */
                {8'h31,8'hb7,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,C,3 */
                {8'h31,8'hc7,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,C,4 */
                {8'h31,8'hd7,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,C,5 */
                {8'h31,8'he7,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,C,6 */
                {8'h31,8'hf7,2'bxx} : dec_alu_shl_adrstage = 1'b1;  /* SHL,C,7 */
                default : dec_alu_shl_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_alu_shl <= 1'b0;
        else if(cpuen) dec_alu_shl <= dec_alu_shl_adrstage;
    end
    output dec_alu_sar;
    reg    dec_alu_sar, dec_alu_sar_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_alu_sar_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h31,8'h0b,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SAR,A,0 */
                {8'h31,8'h1b,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SAR,A,1 */
                {8'h31,8'h2b,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SAR,A,2 */
                {8'h31,8'h3b,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SAR,A,3 */
                {8'h31,8'h4b,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SAR,A,4 */
                {8'h31,8'h5b,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SAR,A,5 */
                {8'h31,8'h6b,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SAR,A,6 */
                {8'h31,8'h7b,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SAR,A,7 */
                {8'h31,8'h0f,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SARW,AX,0 */
                {8'h31,8'h1f,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SARW,AX,1 */
                {8'h31,8'h2f,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SARW,AX,2 */
                {8'h31,8'h3f,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SARW,AX,3 */
                {8'h31,8'h4f,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SARW,AX,4 */
                {8'h31,8'h5f,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SARW,AX,5 */
                {8'h31,8'h6f,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SARW,AX,6 */
                {8'h31,8'h7f,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SARW,AX,7 */
                {8'h31,8'h8f,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SARW,AX,8 */
                {8'h31,8'h9f,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SARW,AX,9 */
                {8'h31,8'haf,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SARW,AX,10 */
                {8'h31,8'hbf,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SARW,AX,11 */
                {8'h31,8'hcf,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SARW,AX,12 */
                {8'h31,8'hdf,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SARW,AX,13 */
                {8'h31,8'hef,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SARW,AX,14 */
                {8'h31,8'hff,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SARW,AX,15 */
                {8'h31,8'h8b,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SAR,A,0 */
                {8'h31,8'h9b,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SAR,A,1 */
                {8'h31,8'hab,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SAR,A,2 */
                {8'h31,8'hbb,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SAR,A,3 */
                {8'h31,8'hcb,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SAR,A,4 */
                {8'h31,8'hdb,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SAR,A,5 */
                {8'h31,8'heb,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SAR,A,6 */
                {8'h31,8'hfb,2'bxx} : dec_alu_sar_adrstage = 1'b1;  /* SAR,A,7 */
                default : dec_alu_sar_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_alu_sar <= 1'b0;
        else if(cpuen) dec_alu_sar <= dec_alu_sar_adrstage;
    end
    output dec_alu_mulu;
    reg    dec_alu_mulu, dec_alu_mulu_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_alu_mulu_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'hd6,8'hxx,2'bxx} : dec_alu_mulu_adrstage = 1'b1;  /* MULU,,X */
                default : dec_alu_mulu_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_alu_mulu <= 1'b0;
        else if(cpuen) dec_alu_mulu <= dec_alu_mulu_adrstage;
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*����ADD,ADDC�Υ��ꥢ�������黻�򣲥���å��ܤ��飱����å��ܤ��ѹ�		*/
/*------------------------------------------------------------------------------*/

    output dec_alu_carry;
    reg    dec_alu_carry, dec_alu_carry_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_alu_carry_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h1c,8'hxx,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,A,#byte */
                {8'h1a,8'hxx,2'bx0} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,saddr,#byte */
                {8'h61,8'h18,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,A,X */
                {8'h61,8'h1a,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,A,C */
                {8'h61,8'h1b,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,A,B */
                {8'h61,8'h1c,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,A,E */
                {8'h61,8'h1d,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,A,D */
                {8'h61,8'h1e,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,A,L */
                {8'h61,8'h1f,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,A,H */
                {8'h61,8'h10,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,X,A */
                {8'h61,8'h11,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,A,A */
                {8'h61,8'h12,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,C,A */
                {8'h61,8'h13,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,B,A */
                {8'h61,8'h14,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,E,A */
                {8'h61,8'h15,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,D,A */
                {8'h61,8'h16,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,L,A */
                {8'h61,8'h17,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,H,A */
                {8'h1b,8'hxx,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,A,saddr */
                {8'h1f,8'hxx,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,A,!addr16 */
                {8'h1d,8'hxx,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,A,[HL] */
                {8'h1e,8'hxx,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,A,[HL+byte] */
                {8'h61,8'h90,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,A,[HL+B] */
                {8'h61,8'h92,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,A,[HL+C] */
                {8'h3c,8'hxx,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,A,#byte */
                {8'h3a,8'hxx,2'bx0} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,saddr,#byte */
                {8'h61,8'h38,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,A,X */
                {8'h61,8'h3a,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,A,C */
                {8'h61,8'h3b,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,A,B */
                {8'h61,8'h3c,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,A,E */
                {8'h61,8'h3d,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,A,D */
                {8'h61,8'h3e,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,A,L */
                {8'h61,8'h3f,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,A,H */
                {8'h61,8'h30,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,X,A */
                {8'h61,8'h31,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,A,A */
                {8'h61,8'h32,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,C,A */
                {8'h61,8'h33,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,B,A */
                {8'h61,8'h34,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,E,A */
                {8'h61,8'h35,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,D,A */
                {8'h61,8'h36,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,L,A */
                {8'h61,8'h37,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,H,A */
                {8'h3b,8'hxx,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,A,saddr */
                {8'h3f,8'hxx,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,A,!addr16 */
                {8'h3d,8'hxx,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,A,[HL] */
                {8'h3e,8'hxx,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,A,[HL+byte] */
                {8'h61,8'hb0,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,A,[HL+B] */
                {8'h61,8'hb2,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,A,[HL+C] */
                {8'h61,8'hfb,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* RORC,A,1 */
                {8'h61,8'hdc,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ROLC,A,1 */
                {8'h61,8'hee,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ROLWC,AX,1 */
                {8'h61,8'hfe,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ROLWC,BC,1 */
                {8'h61,8'h19,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,A,A */
                {8'h61,8'h39,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,A,A */
                {8'h61,8'h91,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,A,[HL+B] */
                {8'h61,8'hb1,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,A,[HL+B] */
                {8'h61,8'h93,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* ADDC,A,[HL+C] */
                {8'h61,8'hb3,2'bxx} : dec_alu_carry_adrstage = 1'b1;  /* SUBC,A,[HL+C] */
                default : dec_alu_carry_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_alu_carry <= 1'b0;
        else if(cpuen) dec_alu_carry <= dec_alu_carry_adrstage;
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*����ž��̿��Ϥ����Ѳ�(MDW�ؽ���+�쥸����)�����Ѳ�				*/
/*------------------------------------------------------------------------------*/

    output [3:0] dec_alu_transout;
    reg    [3:0] dec_alu_transout, dec_alu_transout_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1) begin
            dec_alu_transout_adrstage = 4'h0;
        end else if(ivack == 1'b1) begin
            casex ({stage_adr})  
                {2'b00} : dec_alu_transout_adrstage = 4'hd;  /* Interrupt */
                {2'b01} : dec_alu_transout_adrstage = 4'he;  /* Interrupt */
                default : dec_alu_transout_adrstage = 4'h0;
            endcase
        end else if(skpack == 1'b1) begin
            dec_alu_transout_adrstage = 4'h0;
        end else begin
            if(ID_stage0 == 8'h61) begin
                casex ({ID_stage1,stage_adr})  
                    {8'hd9,2'bxx} : dec_alu_transout_adrstage = 4'h2;  /* MOV,[HL+B],A */
                    {8'hf9,2'bxx} : dec_alu_transout_adrstage = 4'h2;  /* MOV,[HL+C],A */
                    {8'hce,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* MOVS,[HL+byte],X */
                    {8'h8a,2'bxx} : dec_alu_transout_adrstage = 4'h5;  /* XCH,A,C */
                    {8'h8b,2'bxx} : dec_alu_transout_adrstage = 4'h4;  /* XCH,A,B */
                    {8'h8c,2'bxx} : dec_alu_transout_adrstage = 4'h7;  /* XCH,A,E */
                    {8'h8d,2'bxx} : dec_alu_transout_adrstage = 4'h6;  /* XCH,A,D */
                    {8'h8e,2'bxx} : dec_alu_transout_adrstage = 4'h9;  /* XCH,A,L */
                    {8'h8f,2'bxx} : dec_alu_transout_adrstage = 4'h8;  /* XCH,A,H */
                    {8'ha8,2'bx1} : dec_alu_transout_adrstage = 4'h2;  /* XCH,A,saddr */
                    {8'hab,2'bx1} : dec_alu_transout_adrstage = 4'h2;  /* XCH,A,sfr */
                    {8'haa,2'bx1} : dec_alu_transout_adrstage = 4'h2;  /* XCH,A,!addr16 */
                    {8'hae,2'bx1} : dec_alu_transout_adrstage = 4'h2;  /* XCH,A,[DE] */
                    {8'haf,2'bx1} : dec_alu_transout_adrstage = 4'h2;  /* XCH,A,[DE+byte] */
                    {8'hac,2'bx1} : dec_alu_transout_adrstage = 4'h2;  /* XCH,A,[HL] */
                    {8'had,2'bx1} : dec_alu_transout_adrstage = 4'h2;  /* XCH,A,[HL+byte] */
                    {8'hb9,2'bx1} : dec_alu_transout_adrstage = 4'h2;  /* XCH,A,[HL+B] */
                    {8'ha9,2'bx1} : dec_alu_transout_adrstage = 4'h2;  /* XCH,A,[HL+C] */
                    {8'h88,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* XCH,A,X */
                    {8'h98,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* XCH,A,X */
                    {8'h99,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* XCH,A,X */
                    {8'h9a,2'bxx} : dec_alu_transout_adrstage = 4'h5;  /* XCH,A,C */
                    {8'h9b,2'bxx} : dec_alu_transout_adrstage = 4'h4;  /* XCH,A,B */
                    {8'h9c,2'bxx} : dec_alu_transout_adrstage = 4'h7;  /* XCH,A,E */
                    {8'h9d,2'bxx} : dec_alu_transout_adrstage = 4'h6;  /* XCH,A,D */
                    {8'h9e,2'bxx} : dec_alu_transout_adrstage = 4'h9;  /* XCH,A,L */
                    {8'h9f,2'bxx} : dec_alu_transout_adrstage = 4'h8;  /* XCH,A,H */
                    {8'hbb,2'bx1} : dec_alu_transout_adrstage = 4'h2;  /* XCH,A,sfr */
                    {8'hba,2'bx1} : dec_alu_transout_adrstage = 4'h2;  /* XCH,A,!addr16 */
                    {8'hbe,2'bx1} : dec_alu_transout_adrstage = 4'h2;  /* XCH,A,[DE] */
                    {8'hbf,2'bx1} : dec_alu_transout_adrstage = 4'h2;  /* XCH,A,[DE+byte] */
                    {8'hbc,2'bx1} : dec_alu_transout_adrstage = 4'h2;  /* XCH,A,[HL] */
                    {8'hbd,2'bx1} : dec_alu_transout_adrstage = 4'h2;  /* XCH,A,[HL+byte] */
                    {8'h59,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* INC,,[HL+byte] */
                    {8'h69,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* DEC,,[HL+byte] */
                    {8'h79,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* INCW,,[HL+byte] */
                    {8'h89,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* DECW,,[HL+byte] */
                    {8'hca,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALL,,AX */
                    {8'hca,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALL,,AX */
                    {8'hda,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALL,,BC */
                    {8'hda,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALL,,BC */
                    {8'hea,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALL,,DE */
                    {8'hea,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALL,,DE */
                    {8'hfa,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALL,,HL */
                    {8'hfa,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALL,,HL */
                    {8'h84,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[0080h] */
                    {8'h84,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[0080h] */
                    {8'h94,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[0082h] */
                    {8'h94,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[0082h] */
                    {8'ha4,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[0084h] */
                    {8'ha4,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[0084h] */
                    {8'hb4,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[0086h] */
                    {8'hb4,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[0086h] */
                    {8'hc4,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[0088h] */
                    {8'hc4,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[0088h] */
                    {8'hd4,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[008Ah] */
                    {8'hd4,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[008Ah] */
                    {8'he4,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[008Ch] */
                    {8'he4,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[008Ch] */
                    {8'hf4,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[008Eh] */
                    {8'hf4,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[008Eh] */
                    {8'h85,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[0090h] */
                    {8'h85,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[0090h] */
                    {8'h95,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[0092h] */
                    {8'h95,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[0092h] */
                    {8'ha5,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[0094h] */
                    {8'ha5,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[0094h] */
                    {8'hb5,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[0096h] */
                    {8'hb5,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[0096h] */
                    {8'hc5,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[0098h] */
                    {8'hc5,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[0098h] */
                    {8'hd5,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[009Ah] */
                    {8'hd5,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[009Ah] */
                    {8'he5,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[009Ch] */
                    {8'he5,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[009Ch] */
                    {8'hf5,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[009Eh] */
                    {8'hf5,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[009Eh] */
                    {8'h86,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[00A0h] */
                    {8'h86,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[00A0h] */
                    {8'h96,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[00A2h] */
                    {8'h96,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[00A2h] */
                    {8'ha6,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[00A4h] */
                    {8'ha6,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[00A4h] */
                    {8'hb6,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[00A6h] */
                    {8'hb6,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[00A6h] */
                    {8'hc6,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[00A8h] */
                    {8'hc6,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[00A8h] */
                    {8'hd6,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[00AAh] */
                    {8'hd6,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[00AAh] */
                    {8'he6,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[00ACh] */
                    {8'he6,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[00ACh] */
                    {8'hf6,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[00AEh] */
                    {8'hf6,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[00AEh] */
                    {8'h87,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[00B0h] */
                    {8'h87,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[00B0h] */
                    {8'h97,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[00B2h] */
                    {8'h97,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[00B2h] */
                    {8'ha7,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[00B4h] */
                    {8'ha7,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[00B4h] */
                    {8'hb7,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[00B6h] */
                    {8'hb7,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[00B6h] */
                    {8'hc7,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[00B8h] */
                    {8'hc7,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[00B8h] */
                    {8'hd7,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[00BAh] */
                    {8'hd7,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[00BAh] */
                    {8'he7,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[00BCh] */
                    {8'he7,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[00BCh] */
                    {8'hf7,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALLT,,[00BEh] */
                    {8'hf7,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALLT,,[00BEh] */
                    {8'hcc,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* BRK,, */
                    {8'hcc,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* BRK,, */
                    {8'hdd,2'bxx} : dec_alu_transout_adrstage = 4'hf;  /* PUSH,,PSW */
                    {8'ha1,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* SOFT2,,BREAK */
                    {8'ha1,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SOFT2,,BREAK */
                    {8'hb1,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* SOFT3,,BREAK */
                    {8'hb1,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SOFT3,,BREAK */
                    {8'hc1,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* SOFT4,,BREAK */
                    {8'hc1,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SOFT4,,BREAK */
                    default : dec_alu_transout_adrstage = 4'h0;
                endcase
            end else if(ID_stage0 == 8'h71) begin
                casex ({ID_stage1,stage_adr})  
                    {8'h01,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,saddr.0,CY */
                    {8'h11,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,saddr.1,CY */
                    {8'h21,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,saddr.2,CY */
                    {8'h31,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,saddr.3,CY */
                    {8'h41,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,saddr.4,CY */
                    {8'h51,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,saddr.5,CY */
                    {8'h61,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,saddr.6,CY */
                    {8'h71,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,saddr.7,CY */
                    {8'h09,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,sfr.0,CY */
                    {8'h19,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,sfr.1,CY */
                    {8'h29,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,sfr.2,CY */
                    {8'h39,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,sfr.3,CY */
                    {8'h49,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,sfr.4,CY */
                    {8'h59,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,sfr.5,CY */
                    {8'h69,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,sfr.6,CY */
                    {8'h79,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,sfr.7,CY */
                    {8'h81,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,[HL].0,CY */
                    {8'h91,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,[HL].1,CY */
                    {8'ha1,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,[HL].2,CY */
                    {8'hb1,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,[HL].3,CY */
                    {8'hc1,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,[HL].4,CY */
                    {8'hd1,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,[HL].5,CY */
                    {8'he1,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,[HL].6,CY */
                    {8'hf1,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* MOV1,[HL].7,CY */
                    {8'h02,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,saddr.0 */
                    {8'h12,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,saddr.1 */
                    {8'h22,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,saddr.2 */
                    {8'h32,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,saddr.3 */
                    {8'h42,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,saddr.4 */
                    {8'h52,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,saddr.5 */
                    {8'h62,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,saddr.6 */
                    {8'h72,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,saddr.7 */
                    {8'h0a,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,sfr.0 */
                    {8'h1a,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,sfr.1 */
                    {8'h2a,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,sfr.2 */
                    {8'h3a,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,sfr.3 */
                    {8'h4a,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,sfr.4 */
                    {8'h5a,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,sfr.5 */
                    {8'h6a,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,sfr.6 */
                    {8'h7a,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,sfr.7 */
                    {8'h00,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,!addr16.0 */
                    {8'h10,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,!addr16.1 */
                    {8'h20,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,!addr16.2 */
                    {8'h30,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,!addr16.3 */
                    {8'h40,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,!addr16.4 */
                    {8'h50,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,!addr16.5 */
                    {8'h60,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,!addr16.6 */
                    {8'h70,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,!addr16.7 */
                    {8'h82,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,[HL].0 */
                    {8'h92,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,[HL].1 */
                    {8'ha2,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,[HL].2 */
                    {8'hb2,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,[HL].3 */
                    {8'hc2,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,[HL].4 */
                    {8'hd2,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,[HL].5 */
                    {8'he2,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,[HL].6 */
                    {8'hf2,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SET1,,[HL].7 */
                    {8'h03,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,saddr.0 */
                    {8'h13,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,saddr.1 */
                    {8'h23,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,saddr.2 */
                    {8'h33,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,saddr.3 */
                    {8'h43,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,saddr.4 */
                    {8'h53,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,saddr.5 */
                    {8'h63,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,saddr.6 */
                    {8'h73,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,saddr.7 */
                    {8'h0b,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,sfr.0 */
                    {8'h1b,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,sfr.1 */
                    {8'h2b,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,sfr.2 */
                    {8'h3b,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,sfr.3 */
                    {8'h4b,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,sfr.4 */
                    {8'h5b,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,sfr.5 */
                    {8'h6b,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,sfr.6 */
                    {8'h7b,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,sfr.7 */
                    {8'h08,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,!addr16.0 */
                    {8'h18,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,!addr16.1 */
                    {8'h28,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,!addr16.2 */
                    {8'h38,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,!addr16.3 */
                    {8'h48,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,!addr16.4 */
                    {8'h58,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,!addr16.5 */
                    {8'h68,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,!addr16.6 */
                    {8'h78,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,!addr16.7 */
                    {8'h83,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,[HL].0 */
                    {8'h93,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,[HL].1 */
                    {8'ha3,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,[HL].2 */
                    {8'hb3,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,[HL].3 */
                    {8'hc3,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,[HL].4 */
                    {8'hd3,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,[HL].5 */
                    {8'he3,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,[HL].6 */
                    {8'hf3,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CLR1,,[HL].7 */
                    default : dec_alu_transout_adrstage = 4'h0;
                endcase
            end else if(ID_stage0 == 8'h31) begin
                casex ({ID_stage1,stage_adr})  
                    {8'h00,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,saddr.0,$addr8 */
                    {8'h10,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,saddr.1,$addr8 */
                    {8'h20,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,saddr.2,$addr8 */
                    {8'h30,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,saddr.3,$addr8 */
                    {8'h40,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,saddr.4,$addr8 */
                    {8'h50,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,saddr.5,$addr8 */
                    {8'h60,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,saddr.6,$addr8 */
                    {8'h70,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,saddr.7,$addr8 */
                    {8'h80,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,sfr.0,$addr8 */
                    {8'h90,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,sfr.1,$addr8 */
                    {8'ha0,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,sfr.2,$addr8 */
                    {8'hb0,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,sfr.3,$addr8 */
                    {8'hc0,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,sfr.4,$addr8 */
                    {8'hd0,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,sfr.5,$addr8 */
                    {8'he0,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,sfr.6,$addr8 */
                    {8'hf0,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,sfr.7,$addr8 */
                    {8'h81,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,[HL].0,$addr8 */
                    {8'h91,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,[HL].1,$addr8 */
                    {8'ha1,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,[HL].2,$addr8 */
                    {8'hb1,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,[HL].3,$addr8 */
                    {8'hc1,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,[HL].4,$addr8 */
                    {8'hd1,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,[HL].5,$addr8 */
                    {8'he1,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,[HL].6,$addr8 */
                    {8'hf1,2'b10} : dec_alu_transout_adrstage = 4'he;  /* BTCLR,[HL].7,$addr8 */
                    default : dec_alu_transout_adrstage = 4'h0;
                endcase
            end else begin
                casex ({ID_stage0,stage_adr})  
                    {8'h50,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOV,X,#byte */
                    {8'h51,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOV,A,#byte */
                    {8'h52,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOV,C,#byte */
                    {8'h53,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOV,B,#byte */
                    {8'h54,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOV,E,#byte */
                    {8'h55,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOV,D,#byte */
                    {8'h56,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOV,L,#byte */
                    {8'h57,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOV,H,#byte */
                    {8'hcd,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOV,saddr,#byte */
                    {8'hce,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOV,sfr,#byte */
                    {8'hcf,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOV,!addr16,#byte */
                    {8'hca,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOV,[DE+byte],#byte */
                    {8'hcc,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOV,[HL+byte],#byte */
                    {8'h60,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* MOV,A,X */
                    {8'h62,2'bxx} : dec_alu_transout_adrstage = 4'h5;  /* MOV,A,C */
                    {8'h63,2'bxx} : dec_alu_transout_adrstage = 4'h4;  /* MOV,A,B */
                    {8'h64,2'bxx} : dec_alu_transout_adrstage = 4'h7;  /* MOV,A,E */
                    {8'h65,2'bxx} : dec_alu_transout_adrstage = 4'h6;  /* MOV,A,D */
                    {8'h66,2'bxx} : dec_alu_transout_adrstage = 4'h9;  /* MOV,A,L */
                    {8'h67,2'bxx} : dec_alu_transout_adrstage = 4'h8;  /* MOV,A,H */
                    {8'h70,2'bxx} : dec_alu_transout_adrstage = 4'h2;  /* MOV,X,A */
                    {8'h72,2'bxx} : dec_alu_transout_adrstage = 4'h2;  /* MOV,C,A */
                    {8'h73,2'bxx} : dec_alu_transout_adrstage = 4'h2;  /* MOV,B,A */
                    {8'h74,2'bxx} : dec_alu_transout_adrstage = 4'h2;  /* MOV,E,A */
                    {8'h75,2'bxx} : dec_alu_transout_adrstage = 4'h2;  /* MOV,D,A */
                    {8'h76,2'bxx} : dec_alu_transout_adrstage = 4'h2;  /* MOV,L,A */
                    {8'h77,2'bxx} : dec_alu_transout_adrstage = 4'h2;  /* MOV,H,A */
                    {8'h9d,2'bxx} : dec_alu_transout_adrstage = 4'h2;  /* MOV,saddr,A */
                    {8'h9e,2'bxx} : dec_alu_transout_adrstage = 4'h2;  /* MOV,sfr,A */
                    {8'h9f,2'bxx} : dec_alu_transout_adrstage = 4'h2;  /* MOV,!addr16,A */
                    {8'h41,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOV,ES,#byte */
                    {8'h99,2'bxx} : dec_alu_transout_adrstage = 4'h2;  /* MOV,[DE],A */
                    {8'h9a,2'bxx} : dec_alu_transout_adrstage = 4'h2;  /* MOV,[DE+byte],A */
                    {8'h9b,2'bxx} : dec_alu_transout_adrstage = 4'h2;  /* MOV,[HL],A */
                    {8'h9c,2'bxx} : dec_alu_transout_adrstage = 4'h2;  /* MOV,[HL+byte],A */
                    {8'h19,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOV,word[B],#byte */
                    {8'h18,2'bxx} : dec_alu_transout_adrstage = 4'h2;  /* MOV,word[B],A */
                    {8'h38,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOV,word[C],#byte */
                    {8'h28,2'bxx} : dec_alu_transout_adrstage = 4'h2;  /* MOV,word[C],A */
                    {8'h39,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOV,word[BC],#byte */
                    {8'h48,2'bxx} : dec_alu_transout_adrstage = 4'h2;  /* MOV,word[BC],A */
                    {8'hc8,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOV,[SP+byte],#byte */
                    {8'h98,2'bxx} : dec_alu_transout_adrstage = 4'h2;  /* MOV,[SP+byte],A */
                    {8'h08,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* XCH,A,X */
                    {8'h30,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOVW,AX,#word */
                    {8'h32,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOVW,BC,#word */
                    {8'h34,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOVW,DE,#word */
                    {8'h36,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOVW,HL,#word */
                    {8'hc9,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOVW,saddrp,#word */
                    {8'hcb,2'bxx} : dec_alu_transout_adrstage = 4'ha;  /* MOVW,sfrp,#word */
                    {8'hbd,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* MOVW,saddrp,AX */
                    {8'hbe,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* MOVW,sfrp,AX */
                    {8'h13,2'bxx} : dec_alu_transout_adrstage = 4'h5;  /* MOVW,AX,BC */
                    {8'h12,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* MOVW,BC,AX */
                    {8'h15,2'bxx} : dec_alu_transout_adrstage = 4'h7;  /* MOVW,AX,DE */
                    {8'h14,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* MOVW,DE,AX */
                    {8'h17,2'bxx} : dec_alu_transout_adrstage = 4'h9;  /* MOVW,AX,HL */
                    {8'h16,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* MOVW,HL,AX */
                    {8'hbf,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* MOVW,!addr16,AX */
                    {8'hb9,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* MOVW,[DE],AX */
                    {8'hba,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* MOVW,[DE+byte],AX */
                    {8'hbb,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* MOVW,[HL],AX */
                    {8'hbc,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* MOVW,[HL+byte],AX */
                    {8'h58,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* MOVW,word[B],AX */
                    {8'h68,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* MOVW,word[C],AX */
                    {8'h78,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* MOVW,word[BC],AX */
                    {8'hb8,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* MOVW,[SP+byte],AX */
                    {8'h33,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* XCHW,AX,BC */
                    {8'h35,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* XCHW,AX,DE */
                    {8'h37,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* XCHW,AX,HL */
                    {8'he1,2'bxx} : dec_alu_transout_adrstage = 4'h1;  /* ONEB,,A */
                    {8'he0,2'bxx} : dec_alu_transout_adrstage = 4'h1;  /* ONEB,,X */
                    {8'he3,2'bxx} : dec_alu_transout_adrstage = 4'h1;  /* ONEB,,B */
                    {8'he2,2'bxx} : dec_alu_transout_adrstage = 4'h1;  /* ONEB,,C */
                    {8'he4,2'bxx} : dec_alu_transout_adrstage = 4'h1;  /* ONEB,,saddr */
                    {8'he5,2'bxx} : dec_alu_transout_adrstage = 4'h1;  /* ONEB,,!addr16 */
                    {8'he6,2'bxx} : dec_alu_transout_adrstage = 4'h1;  /* ONEW,,AX */
                    {8'he7,2'bxx} : dec_alu_transout_adrstage = 4'h1;  /* ONEW,,BC */
                    {8'h0a,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* ADD,saddr,#byte */
                    {8'h1a,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* ADDC,saddr,#byte */
                    {8'h2a,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SUB,saddr,#byte */
                    {8'h3a,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SUBC,saddr,#byte */
                    {8'h5a,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* AND,saddr,#byte */
                    {8'h6a,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* OR,saddr,#byte */
                    {8'h7a,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* XOR,saddr,#byte */
                    {8'ha4,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* INC,,saddr */
                    {8'ha0,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* INC,,!addr16 */
                    {8'hb4,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* DEC,,saddr */
                    {8'hb0,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* DEC,,!addr16 */
                    {8'ha6,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* INCW,,saddrp */
                    {8'ha2,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* INCW,,!addr16 */
                    {8'hb6,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* DECW,,saddrp */
                    {8'hb2,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* DECW,,!addr16 */
                    {8'hfe,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALL,,$!addr16 */
                    {8'hfe,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALL,,$!addr16 */
                    {8'hfd,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALL,,!addr16 */
                    {8'hfd,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALL,,!addr16 */
                    {8'hfc,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* CALL,,!!addr20 */
                    {8'hfc,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* CALL,,!!addr20 */
                    {8'hff,2'bx0} : dec_alu_transout_adrstage = 4'hd;  /* SOFT,,BREAK */
                    {8'hff,2'bx1} : dec_alu_transout_adrstage = 4'he;  /* SOFT,,BREAK */
                    {8'hc1,2'bxx} : dec_alu_transout_adrstage = 4'h3;  /* PUSH,,AX */
                    {8'hc3,2'bxx} : dec_alu_transout_adrstage = 4'h5;  /* PUSH,,BC */
                    {8'hc5,2'bxx} : dec_alu_transout_adrstage = 4'h7;  /* PUSH,,DE */
                    {8'hc7,2'bxx} : dec_alu_transout_adrstage = 4'h9;  /* PUSH,,HL */
                    default : dec_alu_transout_adrstage = 4'h0;
                endcase
            end
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_alu_transout <= 4'h0;
        else if(cpuen) dec_alu_transout <= dec_alu_transout_adrstage;
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*����ž��̿��Ϥ����Ѳ�(MDR��������+�쥸����)�����Ѳ�				*/
/*------------------------------------------------------------------------------*/
    output dec_alu_transin;
    reg    dec_alu_transin, dec_alu_transin_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1) begin
            dec_alu_transin_adrstage = 1'b0;
        end else if(ivack == 1'b1) begin
            dec_alu_transin_adrstage = 1'b0;
        end else if(skpack == 1'b1) begin
            dec_alu_transin_adrstage = 1'b0;
        end else begin
            if(ID_stage0 == 8'h61) begin
                casex ({ID_stage1,stage_adr})  
                    {8'hc9,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOV,A,[HL+B] */
                    {8'he9,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOV,A,[HL+C] */
                    {8'hb8,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOV,ES,saddr */
                    {8'ha8,2'bx0} : dec_alu_transin_adrstage = 1'b1;  /* XCH,A,saddr */
                    {8'hab,2'bx0} : dec_alu_transin_adrstage = 1'b1;  /* XCH,A,sfr */
                    {8'haa,2'bx0} : dec_alu_transin_adrstage = 1'b1;  /* XCH,A,!addr16 */
                    {8'hae,2'bx0} : dec_alu_transin_adrstage = 1'b1;  /* XCH,A,[DE] */
                    {8'haf,2'bx0} : dec_alu_transin_adrstage = 1'b1;  /* XCH,A,[DE+byte] */
                    {8'hac,2'bx0} : dec_alu_transin_adrstage = 1'b1;  /* XCH,A,[HL] */
                    {8'had,2'bx0} : dec_alu_transin_adrstage = 1'b1;  /* XCH,A,[HL+byte] */
                    {8'hb9,2'bx0} : dec_alu_transin_adrstage = 1'b1;  /* XCH,A,[HL+B] */
                    {8'ha9,2'bx0} : dec_alu_transin_adrstage = 1'b1;  /* XCH,A,[HL+C] */
                    {8'hbb,2'bx0} : dec_alu_transin_adrstage = 1'b1;  /* XCH,A,sfr */
                    {8'hba,2'bx0} : dec_alu_transin_adrstage = 1'b1;  /* XCH,A,!addr16 */
                    {8'hbe,2'bx0} : dec_alu_transin_adrstage = 1'b1;  /* XCH,A,[DE] */
                    {8'hbf,2'bx0} : dec_alu_transin_adrstage = 1'b1;  /* XCH,A,[DE+byte] */
                    {8'hbc,2'bx0} : dec_alu_transin_adrstage = 1'b1;  /* XCH,A,[HL] */
                    {8'hbd,2'bx0} : dec_alu_transin_adrstage = 1'b1;  /* XCH,A,[HL+byte] */
                    default : dec_alu_transin_adrstage = 1'b0;
                endcase
            end else begin
                casex ({ID_stage0,stage_adr})  
                    {8'h8d,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOV,A,saddr */
                    {8'h8e,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOV,A,sfr */
                    {8'h8f,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOV,A,!addr16 */
                    {8'h89,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOV,A,[DE] */
                    {8'h8a,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOV,A,[DE+byte] */
                    {8'h8b,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOV,A,[HL] */
                    {8'h8c,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOV,A,[HL+byte] */
                    {8'h09,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOV,A,word[B] */
                    {8'h29,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOV,A,word[C] */
                    {8'h49,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOV,A,word[BC] */
                    {8'h88,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOV,A,[SP+byte] */
                    {8'he8,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOV,B,saddr */
                    {8'he9,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOV,B,!addr16 */
                    {8'hf8,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOV,C,saddr */
                    {8'hf9,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOV,C,!addr16 */
                    {8'hd8,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOV,X,saddr */
                    {8'hd9,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOV,X,!addr16 */
                    {8'had,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOVW,AX,saddrp */
                    {8'hae,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOVW,AX,sfrp */
                    {8'haf,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOVW,AX,!addr16 */
                    {8'ha9,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOVW,AX,[DE] */
                    {8'haa,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOVW,AX,[DE+byte] */
                    {8'hab,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOVW,AX,[HL] */
                    {8'hac,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOVW,AX,[HL+byte] */
                    {8'h59,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOVW,AX,word[B] */
                    {8'h69,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOVW,AX,word[C] */
                    {8'h79,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOVW,AX,word[BC] */
                    {8'ha8,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOVW,AX,[SP+byte] */
                    {8'hda,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOVW,BC,saddrp */
                    {8'hdb,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOVW,BC,!addr16 */
                    {8'hea,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOVW,DE,saddrp */
                    {8'heb,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOVW,DE,!addr16 */
                    {8'hfa,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOVW,HL,saddrp */
                    {8'hfb,2'bxx} : dec_alu_transin_adrstage = 1'b1;  /* MOVW,HL,!addr16 */
                    default : dec_alu_transin_adrstage = 1'b0;
                endcase
            end
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_alu_transin <= 1'b0;
        else if(cpuen) dec_alu_transin <= dec_alu_transin_adrstage;
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�������ե�̿��Ϥ����Ѳ�(MDW�ؽ���+�쥸����) �����Ѳ�				*/
/*------------------------------------------------------------------------------*/

    output [4:0] dec_alu_bitsh ;
    reg    [4:0] dec_alu_bitsh ,dec_alu_bitsh_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1) begin
            dec_alu_bitsh_adrstage = 5'h0;
        end else if(ivack == 1'b1) begin
            dec_alu_bitsh_adrstage = 5'h0;
        end else if(skpack == 1'b1) begin
            dec_alu_bitsh_adrstage = 5'h0;
        end else begin
            if(ID_stage0 == 8'h61) begin                               /* ROR, ROL, RORC, ROLC, ROLWC  */
                casex ({ID_stage1,stage_adr})  
                    {8'hdb,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* ROR,A,1 */
                    {8'heb,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* ROL,A,1 */
                    {8'hfb,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* RORC,A,1 */
                    {8'hdc,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* ROLC,A,1 */
                    {8'hee,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* ROLWC,AX,1 */
                    {8'hfe,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* ROLWC,BC,1 */
                    default : dec_alu_bitsh_adrstage = 5'h0;
                endcase
            end else if(ID_stage0 == 8'h71) begin			/* MOV1, AND1, OR1, XOR1, SET1, CLR1, NOT1 */
                casex ({ID_stage1,stage_adr})  
                    {8'h04,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,saddr.0 */
                    {8'h14,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,saddr.1 */
                    {8'h24,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,saddr.2 */
                    {8'h34,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,saddr.3 */
                    {8'h44,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,saddr.4 */
                    {8'h54,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,saddr.5 */
                    {8'h64,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,saddr.6 */
                    {8'h74,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,saddr.7 */
                    {8'h0c,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,sfr.0 */
                    {8'h1c,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,sfr.1 */
                    {8'h2c,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,sfr.2 */
                    {8'h3c,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,sfr.3 */
                    {8'h4c,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,sfr.4 */
                    {8'h5c,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,sfr.5 */
                    {8'h6c,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,sfr.6 */
                    {8'h7c,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,sfr.7 */
                    {8'h8c,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* MOV1,CY,A.0 */
                    {8'h9c,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* MOV1,CY,A.1 */
                    {8'hac,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* MOV1,CY,A.2 */
                    {8'hbc,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* MOV1,CY,A.3 */
                    {8'hcc,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* MOV1,CY,A.4 */
                    {8'hdc,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* MOV1,CY,A.5 */
                    {8'hec,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* MOV1,CY,A.6 */
                    {8'hfc,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* MOV1,CY,A.7 */
                    {8'h84,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,[HL].0 */
                    {8'h94,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,[HL].1 */
                    {8'ha4,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,[HL].2 */
                    {8'hb4,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,[HL].3 */
                    {8'hc4,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,[HL].4 */
                    {8'hd4,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,[HL].5 */
                    {8'he4,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,[HL].6 */
                    {8'hf4,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* MOV1,CY,[HL].7 */
                    {8'h01,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,saddr.0,CY */
                    {8'h11,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,saddr.1,CY */
                    {8'h21,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,saddr.2,CY */
                    {8'h31,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,saddr.3,CY */
                    {8'h41,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,saddr.4,CY */
                    {8'h51,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,saddr.5,CY */
                    {8'h61,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,saddr.6,CY */
                    {8'h71,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,saddr.7,CY */
                    {8'h09,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,sfr.0,CY */
                    {8'h19,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,sfr.1,CY */
                    {8'h29,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,sfr.2,CY */
                    {8'h39,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,sfr.3,CY */
                    {8'h49,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,sfr.4,CY */
                    {8'h59,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,sfr.5,CY */
                    {8'h69,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,sfr.6,CY */
                    {8'h79,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,sfr.7,CY */
                    {8'h89,2'bxx} : dec_alu_bitsh_adrstage = 5'hf;   /* MOV1,A.0,CY */
                    {8'h99,2'bxx} : dec_alu_bitsh_adrstage = 5'hf;   /* MOV1,A.1,CY */
                    {8'ha9,2'bxx} : dec_alu_bitsh_adrstage = 5'hf;   /* MOV1,A.2,CY */
                    {8'hb9,2'bxx} : dec_alu_bitsh_adrstage = 5'hf;   /* MOV1,A.3,CY */
                    {8'hc9,2'bxx} : dec_alu_bitsh_adrstage = 5'hf;   /* MOV1,A.4,CY */
                    {8'hd9,2'bxx} : dec_alu_bitsh_adrstage = 5'hf;   /* MOV1,A.5,CY */
                    {8'he9,2'bxx} : dec_alu_bitsh_adrstage = 5'hf;   /* MOV1,A.6,CY */
                    {8'hf9,2'bxx} : dec_alu_bitsh_adrstage = 5'hf;   /* MOV1,A.7,CY */
                    {8'h81,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,[HL].0,CY */
                    {8'h91,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,[HL].1,CY */
                    {8'ha1,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,[HL].2,CY */
                    {8'hb1,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,[HL].3,CY */
                    {8'hc1,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,[HL].4,CY */
                    {8'hd1,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,[HL].5,CY */
                    {8'he1,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,[HL].6,CY */
                    {8'hf1,2'bx0} : dec_alu_bitsh_adrstage = 5'he;   /* MOV1,[HL].7,CY */
                    {8'h05,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,saddr.0 */
                    {8'h15,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,saddr.1 */
                    {8'h25,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,saddr.2 */
                    {8'h35,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,saddr.3 */
                    {8'h45,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,saddr.4 */
                    {8'h55,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,saddr.5 */
                    {8'h65,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,saddr.6 */
                    {8'h75,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,saddr.7 */
                    {8'h0d,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,sfr.0 */
                    {8'h1d,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,sfr.1 */
                    {8'h2d,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,sfr.2 */
                    {8'h3d,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,sfr.3 */
                    {8'h4d,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,sfr.4 */
                    {8'h5d,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,sfr.5 */
                    {8'h6d,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,sfr.6 */
                    {8'h7d,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,sfr.7 */
                    {8'h8d,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* AND1,CY,A.0 */
                    {8'h9d,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* AND1,CY,A.1 */
                    {8'had,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* AND1,CY,A.2 */
                    {8'hbd,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* AND1,CY,A.3 */
                    {8'hcd,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* AND1,CY,A.4 */
                    {8'hdd,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* AND1,CY,A.5 */
                    {8'hed,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* AND1,CY,A.6 */
                    {8'hfd,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* AND1,CY,A.7 */
                    {8'h85,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,[HL].0 */
                    {8'h95,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,[HL].1 */
                    {8'ha5,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,[HL].2 */
                    {8'hb5,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,[HL].3 */
                    {8'hc5,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,[HL].4 */
                    {8'hd5,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,[HL].5 */
                    {8'he5,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,[HL].6 */
                    {8'hf5,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* AND1,CY,[HL].7 */
                    {8'h06,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,saddr.0 */
                    {8'h16,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,saddr.1 */
                    {8'h26,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,saddr.2 */
                    {8'h36,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,saddr.3 */
                    {8'h46,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,saddr.4 */
                    {8'h56,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,saddr.5 */
                    {8'h66,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,saddr.6 */
                    {8'h76,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,saddr.7 */
                    {8'h0e,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,sfr.0 */
                    {8'h1e,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,sfr.1 */
                    {8'h2e,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,sfr.2 */
                    {8'h3e,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,sfr.3 */
                    {8'h4e,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,sfr.4 */
                    {8'h5e,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,sfr.5 */
                    {8'h6e,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,sfr.6 */
                    {8'h7e,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,sfr.7 */
                    {8'h8e,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* OR1,CY,A.0 */
                    {8'h9e,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* OR1,CY,A.1 */
                    {8'hae,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* OR1,CY,A.2 */
                    {8'hbe,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* OR1,CY,A.3 */
                    {8'hce,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* OR1,CY,A.4 */
                    {8'hde,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* OR1,CY,A.5 */
                    {8'hee,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* OR1,CY,A.6 */
                    {8'hfe,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* OR1,CY,A.7 */
                    {8'h86,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,[HL].0 */
                    {8'h96,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,[HL].1 */
                    {8'ha6,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,[HL].2 */
                    {8'hb6,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,[HL].3 */
                    {8'hc6,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,[HL].4 */
                    {8'hd6,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,[HL].5 */
                    {8'he6,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,[HL].6 */
                    {8'hf6,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* OR1,CY,[HL].7 */
                    {8'h07,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,saddr.0 */
                    {8'h17,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,saddr.1 */
                    {8'h27,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,saddr.2 */
                    {8'h37,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,saddr.3 */
                    {8'h47,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,saddr.4 */
                    {8'h57,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,saddr.5 */
                    {8'h67,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,saddr.6 */
                    {8'h77,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,saddr.7 */
                    {8'h0f,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,sfr.0 */
                    {8'h1f,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,sfr.1 */
                    {8'h2f,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,sfr.2 */
                    {8'h3f,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,sfr.3 */
                    {8'h4f,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,sfr.4 */
                    {8'h5f,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,sfr.5 */
                    {8'h6f,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,sfr.6 */
                    {8'h7f,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,sfr.7 */
                    {8'h8f,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* XOR1,CY,A.0 */
                    {8'h9f,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* XOR1,CY,A.1 */
                    {8'haf,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* XOR1,CY,A.2 */
                    {8'hbf,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* XOR1,CY,A.3 */
                    {8'hcf,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* XOR1,CY,A.4 */
                    {8'hdf,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* XOR1,CY,A.5 */
                    {8'hef,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* XOR1,CY,A.6 */
                    {8'hff,2'bxx} : dec_alu_bitsh_adrstage = 5'h9;  /* XOR1,CY,A.7 */
                    {8'h87,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,[HL].0 */
                    {8'h97,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,[HL].1 */
                    {8'ha7,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,[HL].2 */
                    {8'hb7,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,[HL].3 */
                    {8'hc7,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,[HL].4 */
                    {8'hd7,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,[HL].5 */
                    {8'he7,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,[HL].6 */
                    {8'hf7,2'bxx} : dec_alu_bitsh_adrstage = 5'h8;  /* XOR1,CY,[HL].7 */
                    {8'h02,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,saddr.0 */
                    {8'h12,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,saddr.1 */
                    {8'h22,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,saddr.2 */
                    {8'h32,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,saddr.3 */
                    {8'h42,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,saddr.4 */
                    {8'h52,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,saddr.5 */
                    {8'h62,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,saddr.6 */
                    {8'h72,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,saddr.7 */
                    {8'h0a,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,sfr.0 */
                    {8'h1a,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,sfr.1 */
                    {8'h2a,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,sfr.2 */
                    {8'h3a,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,sfr.3 */
                    {8'h4a,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,sfr.4 */
                    {8'h5a,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,sfr.5 */
                    {8'h6a,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,sfr.6 */
                    {8'h7a,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,sfr.7 */
                    {8'h8a,2'bxx} : dec_alu_bitsh_adrstage = 5'h1d;  /* SET1,,A.0 */
                    {8'h9a,2'bxx} : dec_alu_bitsh_adrstage = 5'h1d;  /* SET1,,A.1 */
                    {8'haa,2'bxx} : dec_alu_bitsh_adrstage = 5'h1d;  /* SET1,,A.2 */
                    {8'hba,2'bxx} : dec_alu_bitsh_adrstage = 5'h1d;  /* SET1,,A.3 */
                    {8'hca,2'bxx} : dec_alu_bitsh_adrstage = 5'h1d;  /* SET1,,A.4 */
                    {8'hda,2'bxx} : dec_alu_bitsh_adrstage = 5'h1d;  /* SET1,,A.5 */
                    {8'hea,2'bxx} : dec_alu_bitsh_adrstage = 5'h1d;  /* SET1,,A.6 */
                    {8'hfa,2'bxx} : dec_alu_bitsh_adrstage = 5'h1d;  /* SET1,,A.7 */
                    {8'h00,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,!addr16.0 */
                    {8'h10,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,!addr16.1 */
                    {8'h20,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,!addr16.2 */
                    {8'h30,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,!addr16.3 */
                    {8'h40,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,!addr16.4 */
                    {8'h50,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,!addr16.5 */
                    {8'h60,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,!addr16.6 */
                    {8'h70,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,!addr16.7 */
                    {8'h82,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,[HL].0 */
                    {8'h92,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,[HL].1 */
                    {8'ha2,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,[HL].2 */
                    {8'hb2,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,[HL].3 */
                    {8'hc2,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,[HL].4 */
                    {8'hd2,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,[HL].5 */
                    {8'he2,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,[HL].6 */
                    {8'hf2,2'bx0} : dec_alu_bitsh_adrstage = 5'hd;  /* SET1,,[HL].7 */
                    {8'h03,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,saddr.0 */
                    {8'h13,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,saddr.1 */
                    {8'h23,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,saddr.2 */
                    {8'h33,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,saddr.3 */
                    {8'h43,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,saddr.4 */
                    {8'h53,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,saddr.5 */
                    {8'h63,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,saddr.6 */
                    {8'h73,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,saddr.7 */
                    {8'h0b,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,sfr.0 */
                    {8'h1b,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,sfr.1 */
                    {8'h2b,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,sfr.2 */
                    {8'h3b,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,sfr.3 */
                    {8'h4b,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,sfr.4 */
                    {8'h5b,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,sfr.5 */
                    {8'h6b,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,sfr.6 */
                    {8'h7b,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,sfr.7 */
                    {8'h8b,2'bxx} : dec_alu_bitsh_adrstage = 5'h1c;  /* CLR1,,A.0 */
                    {8'h9b,2'bxx} : dec_alu_bitsh_adrstage = 5'h1c;  /* CLR1,,A.1 */
                    {8'hab,2'bxx} : dec_alu_bitsh_adrstage = 5'h1c;  /* CLR1,,A.2 */
                    {8'hbb,2'bxx} : dec_alu_bitsh_adrstage = 5'h1c;  /* CLR1,,A.3 */
                    {8'hcb,2'bxx} : dec_alu_bitsh_adrstage = 5'h1c;  /* CLR1,,A.4 */
                    {8'hdb,2'bxx} : dec_alu_bitsh_adrstage = 5'h1c;  /* CLR1,,A.5 */
                    {8'heb,2'bxx} : dec_alu_bitsh_adrstage = 5'h1c;  /* CLR1,,A.6 */
                    {8'hfb,2'bxx} : dec_alu_bitsh_adrstage = 5'h1c;  /* CLR1,,A.7 */
                    {8'h08,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,!addr16.0 */
                    {8'h18,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,!addr16.1 */
                    {8'h28,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,!addr16.2 */
                    {8'h38,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,!addr16.3 */
                    {8'h48,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,!addr16.4 */
                    {8'h58,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,!addr16.5 */
                    {8'h68,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,!addr16.6 */
                    {8'h78,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,!addr16.7 */
                    {8'h83,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,[HL].0 */
                    {8'h93,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,[HL].1 */
                    {8'ha3,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,[HL].2 */
                    {8'hb3,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,[HL].3 */
                    {8'hc3,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,[HL].4 */
                    {8'hd3,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,[HL].5 */
                    {8'he3,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,[HL].6 */
                    {8'hf3,2'bx0} : dec_alu_bitsh_adrstage = 5'hc;  /* CLR1,,[HL].7 */
                    {8'h80,2'bxx} : dec_alu_bitsh_adrstage = 5'h1;   /* SET1,,CY */
                    {8'h88,2'bxx} : dec_alu_bitsh_adrstage = 5'h1;   /* CLR1,,CY */
                    {8'hc0,2'bxx} : dec_alu_bitsh_adrstage = 5'h11;  /* NOT1,,CY */
                    {8'h90,2'bxx} : dec_alu_bitsh_adrstage = 5'h1;   /* SET1,,CY */
                    {8'ha0,2'bxx} : dec_alu_bitsh_adrstage = 5'h1;   /* SET1,,CY */
                    {8'hb0,2'bxx} : dec_alu_bitsh_adrstage = 5'h1;   /* SET1,,CY */
                    {8'hd0,2'bxx} : dec_alu_bitsh_adrstage = 5'h11;  /* NOT1,,CY */
                    {8'he0,2'bxx} : dec_alu_bitsh_adrstage = 5'h11;  /* NOT1,,CY */
                    {8'hf0,2'bxx} : dec_alu_bitsh_adrstage = 5'h11;  /* NOT1,,CY */
                    {8'h98,2'bxx} : dec_alu_bitsh_adrstage = 5'h1;   /* CLR1,,CY */
                    {8'ha8,2'bxx} : dec_alu_bitsh_adrstage = 5'h1;   /* CLR1,,CY */
                    {8'hb8,2'bxx} : dec_alu_bitsh_adrstage = 5'h1;   /* CLR1,,CY */
                    {8'hc8,2'bxx} : dec_alu_bitsh_adrstage = 5'h11;  /* NOT1,,CY */
                    {8'hd8,2'bxx} : dec_alu_bitsh_adrstage = 5'h11;  /* NOT1,,CY */
                    {8'he8,2'bxx} : dec_alu_bitsh_adrstage = 5'h11;  /* NOT1,,CY */
                    {8'hf8,2'bxx} : dec_alu_bitsh_adrstage = 5'h11;  /* NOT1,,CY */
                     default : dec_alu_bitsh_adrstage = 5'h0;
                endcase
            end else if(ID_stage0 == 8'h31) begin                      /* SHR, SHRW, SHL, SHLW, SAR, SARW, BT, BF, BTCLR */
                casex ({ID_stage1,stage_adr})  
                    {8'h0a,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHR,A,0 */
                    {8'h1a,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHR,A,1 */
                    {8'h2a,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHR,A,2 */
                    {8'h3a,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHR,A,3 */
                    {8'h4a,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHR,A,4 */
                    {8'h5a,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHR,A,5 */
                    {8'h6a,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHR,A,6 */
                    {8'h7a,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHR,A,7 */
                    {8'h0e,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHRW,AX,0 */
                    {8'h1e,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHRW,AX,1 */
                    {8'h2e,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHRW,AX,2 */
                    {8'h3e,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHRW,AX,3 */
                    {8'h4e,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHRW,AX,4 */
                    {8'h5e,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHRW,AX,5 */
                    {8'h6e,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHRW,AX,6 */
                    {8'h7e,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHRW,AX,7 */
                    {8'h8e,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHRW,AX,8 */
                    {8'h9e,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHRW,AX,9 */
                    {8'hae,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHRW,AX,10 */
                    {8'hbe,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHRW,AX,11 */
                    {8'hce,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHRW,AX,12 */
                    {8'hde,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHRW,AX,13 */
                    {8'hee,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHRW,AX,14 */
                    {8'hfe,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHRW,AX,15 */
                    {8'h09,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHL,A,0 */
                    {8'h19,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHL,A,1 */
                    {8'h29,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHL,A,2 */
                    {8'h39,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHL,A,3 */
                    {8'h49,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHL,A,4 */
                    {8'h59,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHL,A,5 */
                    {8'h69,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHL,A,6 */
                    {8'h79,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHL,A,7 */
                    {8'h08,2'bxx} : dec_alu_bitsh_adrstage = 5'h4;  /* SHL,B,0 */
                    {8'h18,2'bxx} : dec_alu_bitsh_adrstage = 5'h4;  /* SHL,B,1 */
                    {8'h28,2'bxx} : dec_alu_bitsh_adrstage = 5'h4;  /* SHL,B,2 */
                    {8'h38,2'bxx} : dec_alu_bitsh_adrstage = 5'h4;  /* SHL,B,3 */
                    {8'h48,2'bxx} : dec_alu_bitsh_adrstage = 5'h4;  /* SHL,B,4 */
                    {8'h58,2'bxx} : dec_alu_bitsh_adrstage = 5'h4;  /* SHL,B,5 */
                    {8'h68,2'bxx} : dec_alu_bitsh_adrstage = 5'h4;  /* SHL,B,6 */
                    {8'h78,2'bxx} : dec_alu_bitsh_adrstage = 5'h4;  /* SHL,B,7 */
                    {8'h07,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHL,C,0 */
                    {8'h17,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHL,C,1 */
                    {8'h27,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHL,C,2 */
                    {8'h37,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHL,C,3 */
                    {8'h47,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHL,C,4 */
                    {8'h57,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHL,C,5 */
                    {8'h67,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHL,C,6 */
                    {8'h77,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHL,C,7 */
                    {8'h0d,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHLW,AX,0 */
                    {8'h1d,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHLW,AX,1 */
                    {8'h2d,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHLW,AX,2 */
                    {8'h3d,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHLW,AX,3 */
                    {8'h4d,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHLW,AX,4 */
                    {8'h5d,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHLW,AX,5 */
                    {8'h6d,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHLW,AX,6 */
                    {8'h7d,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHLW,AX,7 */
                    {8'h8d,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHLW,AX,8 */
                    {8'h9d,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHLW,AX,9 */
                    {8'had,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHLW,AX,10 */
                    {8'hbd,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHLW,AX,11 */
                    {8'hcd,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHLW,AX,12 */
                    {8'hdd,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHLW,AX,13 */
                    {8'hed,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHLW,AX,14 */
                    {8'hfd,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SHLW,AX,15 */
                    {8'h0c,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHLW,BC,0 */
                    {8'h1c,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHLW,BC,1 */
                    {8'h2c,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHLW,BC,2 */
                    {8'h3c,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHLW,BC,3 */
                    {8'h4c,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHLW,BC,4 */
                    {8'h5c,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHLW,BC,5 */
                    {8'h6c,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHLW,BC,6 */
                    {8'h7c,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHLW,BC,7 */
                    {8'h8c,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHLW,BC,8 */
                    {8'h9c,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHLW,BC,9 */
                    {8'hac,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHLW,BC,10 */
                    {8'hbc,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHLW,BC,11 */
                    {8'hcc,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHLW,BC,12 */
                    {8'hdc,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHLW,BC,13 */
                    {8'hec,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHLW,BC,14 */
                    {8'hfc,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHLW,BC,15 */
                    {8'h0b,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SAR,A,0 */
                    {8'h1b,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SAR,A,1 */
                    {8'h2b,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SAR,A,2 */
                    {8'h3b,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SAR,A,3 */
                    {8'h4b,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SAR,A,4 */
                    {8'h5b,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SAR,A,5 */
                    {8'h6b,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SAR,A,6 */
                    {8'h7b,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SAR,A,7 */
                    {8'h0f,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SARW,AX,0 */
                    {8'h1f,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SARW,AX,1 */
                    {8'h2f,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SARW,AX,2 */
                    {8'h3f,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SARW,AX,3 */
                    {8'h4f,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SARW,AX,4 */
                    {8'h5f,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SARW,AX,5 */
                    {8'h6f,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SARW,AX,6 */
                    {8'h7f,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SARW,AX,7 */
                    {8'h8f,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SARW,AX,8 */
                    {8'h9f,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SARW,AX,9 */
                    {8'haf,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SARW,AX,10 */
                    {8'hbf,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SARW,AX,11 */
                    {8'hcf,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SARW,AX,12 */
                    {8'hdf,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SARW,AX,13 */
                    {8'hef,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SARW,AX,14 */
                    {8'hff,2'bxx} : dec_alu_bitsh_adrstage = 5'h3;  /* SARW,AX,15 */
                    {8'h02,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,saddr.0,$addr8 */
                    {8'h12,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,saddr.1,$addr8 */
                    {8'h22,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,saddr.2,$addr8 */
                    {8'h32,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,saddr.3,$addr8 */
                    {8'h42,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,saddr.4,$addr8 */
                    {8'h52,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,saddr.5,$addr8 */
                    {8'h62,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,saddr.6,$addr8 */
                    {8'h72,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,saddr.7,$addr8 */
                    {8'h82,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,sfr.0,$addr8 */
                    {8'h92,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,sfr.1,$addr8 */
                    {8'ha2,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,sfr.2,$addr8 */
                    {8'hb2,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,sfr.3,$addr8 */
                    {8'hc2,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,sfr.4,$addr8 */
                    {8'hd2,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,sfr.5,$addr8 */
                    {8'he2,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,sfr.6,$addr8 */
                    {8'hf2,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,sfr.7,$addr8 */
                    {8'h03,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BT,A.0,$addr8 */
                    {8'h13,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BT,A.1,$addr8 */
                    {8'h23,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BT,A.2,$addr8 */
                    {8'h33,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BT,A.3,$addr8 */
                    {8'h43,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BT,A.4,$addr8 */
                    {8'h53,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BT,A.5,$addr8 */
                    {8'h63,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BT,A.6,$addr8 */
                    {8'h73,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BT,A.7,$addr8 */
                    {8'h83,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,[HL].0,$addr8 */
                    {8'h93,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,[HL].1,$addr8 */
                    {8'ha3,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,[HL].2,$addr8 */
                    {8'hb3,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,[HL].3,$addr8 */
                    {8'hc3,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,[HL].4,$addr8 */
                    {8'hd3,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,[HL].5,$addr8 */
                    {8'he3,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,[HL].6,$addr8 */
                    {8'hf3,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BT,[HL].7,$addr8 */
                    {8'h04,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,saddr.0,$addr8 */
                    {8'h14,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,saddr.1,$addr8 */
                    {8'h24,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,saddr.2,$addr8 */
                    {8'h34,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,saddr.3,$addr8 */
                    {8'h44,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,saddr.4,$addr8 */
                    {8'h54,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,saddr.5,$addr8 */
                    {8'h64,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,saddr.6,$addr8 */
                    {8'h74,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,saddr.7,$addr8 */
                    {8'h84,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,sfr.0,$addr8 */
                    {8'h94,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,sfr.1,$addr8 */
                    {8'ha4,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,sfr.2,$addr8 */
                    {8'hb4,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,sfr.3,$addr8 */
                    {8'hc4,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,sfr.4,$addr8 */
                    {8'hd4,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,sfr.5,$addr8 */
                    {8'he4,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,sfr.6,$addr8 */
                    {8'hf4,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,sfr.7,$addr8 */
                    {8'h05,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BF,A.0,$addr8 */
                    {8'h15,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BF,A.1,$addr8 */
                    {8'h25,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BF,A.2,$addr8 */
                    {8'h35,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BF,A.3,$addr8 */
                    {8'h45,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BF,A.4,$addr8 */
                    {8'h55,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BF,A.5,$addr8 */
                    {8'h65,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BF,A.6,$addr8 */
                    {8'h75,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BF,A.7,$addr8 */
                    {8'h85,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,[HL].0,$addr8 */
                    {8'h95,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,[HL].1,$addr8 */
                    {8'ha5,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,[HL].2,$addr8 */
                    {8'hb5,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,[HL].3,$addr8 */
                    {8'hc5,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,[HL].4,$addr8 */
                    {8'hd5,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,[HL].5,$addr8 */
                    {8'he5,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,[HL].6,$addr8 */
                    {8'hf5,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BF,[HL].7,$addr8 */
                    {8'h00,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,saddr.0,$addr8 */
                    {8'h00,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,saddr.0,$addr8 */
                    {8'h10,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,saddr.1,$addr8 */
                    {8'h10,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,saddr.1,$addr8 */
                    {8'h20,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,saddr.2,$addr8 */
                    {8'h20,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,saddr.2,$addr8 */
                    {8'h30,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,saddr.3,$addr8 */
                    {8'h30,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,saddr.3,$addr8 */
                    {8'h40,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,saddr.4,$addr8 */
                    {8'h40,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,saddr.4,$addr8 */
                    {8'h50,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,saddr.5,$addr8 */
                    {8'h50,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,saddr.5,$addr8 */
                    {8'h60,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,saddr.6,$addr8 */
                    {8'h60,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,saddr.6,$addr8 */
                    {8'h70,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,saddr.7,$addr8 */
                    {8'h70,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,saddr.7,$addr8 */
                    {8'h80,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,sfr.0,$addr8 */
                    {8'h80,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,sfr.0,$addr8 */
                    {8'h90,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,sfr.1,$addr8 */
                    {8'h90,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,sfr.1,$addr8 */
                    {8'ha0,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,sfr.2,$addr8 */
                    {8'ha0,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,sfr.2,$addr8 */
                    {8'hb0,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,sfr.3,$addr8 */
                    {8'hb0,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,sfr.3,$addr8 */
                    {8'hc0,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,sfr.4,$addr8 */
                    {8'hc0,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,sfr.4,$addr8 */
                    {8'hd0,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,sfr.5,$addr8 */
                    {8'hd0,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,sfr.5,$addr8 */
                    {8'he0,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,sfr.6,$addr8 */
                    {8'he0,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,sfr.6,$addr8 */
                    {8'hf0,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,sfr.7,$addr8 */
                    {8'hf0,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,sfr.7,$addr8 */
                    {8'h01,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BTCLR,A.0,$addr8 */
                    {8'h01,2'b10} : dec_alu_bitsh_adrstage = 5'h1c;  /* BTCLR,A.0,$addr8 */
                    {8'h11,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BTCLR,A.1,$addr8 */
                    {8'h11,2'b10} : dec_alu_bitsh_adrstage = 5'h1c;  /* BTCLR,A.1,$addr8 */
                    {8'h21,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BTCLR,A.2,$addr8 */
                    {8'h21,2'b10} : dec_alu_bitsh_adrstage = 5'h1c;  /* BTCLR,A.2,$addr8 */
                    {8'h31,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BTCLR,A.3,$addr8 */
                    {8'h31,2'b10} : dec_alu_bitsh_adrstage = 5'h1c;  /* BTCLR,A.3,$addr8 */
                    {8'h41,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BTCLR,A.4,$addr8 */
                    {8'h41,2'b10} : dec_alu_bitsh_adrstage = 5'h1c;  /* BTCLR,A.4,$addr8 */
                    {8'h51,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BTCLR,A.5,$addr8 */
                    {8'h51,2'b10} : dec_alu_bitsh_adrstage = 5'h1c;  /* BTCLR,A.5,$addr8 */
                    {8'h61,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BTCLR,A.6,$addr8 */
                    {8'h61,2'b10} : dec_alu_bitsh_adrstage = 5'h1c;  /* BTCLR,A.6,$addr8 */
                    {8'h71,2'b00} : dec_alu_bitsh_adrstage = 5'h19;  /* BTCLR,A.7,$addr8 */
                    {8'h71,2'b10} : dec_alu_bitsh_adrstage = 5'h1c;  /* BTCLR,A.7,$addr8 */
                    {8'h81,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,[HL].0,$addr8 */
                    {8'h81,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,[HL].0,$addr8 */
                    {8'h91,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,[HL].1,$addr8 */
                    {8'h91,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,[HL].1,$addr8 */
                    {8'ha1,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,[HL].2,$addr8 */
                    {8'ha1,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,[HL].2,$addr8 */
                    {8'hb1,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,[HL].3,$addr8 */
                    {8'hb1,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,[HL].3,$addr8 */
                    {8'hc1,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,[HL].4,$addr8 */
                    {8'hc1,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,[HL].4,$addr8 */
                    {8'hd1,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,[HL].5,$addr8 */
                    {8'hd1,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,[HL].5,$addr8 */
                    {8'he1,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,[HL].6,$addr8 */
                    {8'he1,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,[HL].6,$addr8 */
                    {8'hf1,2'b00} : dec_alu_bitsh_adrstage = 5'h18;  /* BTCLR,[HL].7,$addr8 */
                    {8'hf1,2'b01} : dec_alu_bitsh_adrstage = 5'hc;  /* BTCLR,[HL].7,$addr8 */
                    {8'h8a,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHR,A,0 */
                    {8'h9a,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHR,A,1 */
                    {8'haa,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHR,A,2 */
                    {8'hba,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHR,A,3 */
                    {8'hca,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHR,A,4 */
                    {8'hda,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHR,A,5 */
                    {8'hea,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHR,A,6 */
                    {8'hfa,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHR,A,7 */
                    {8'h89,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHL,A,0 */
                    {8'h99,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHL,A,1 */
                    {8'ha9,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHL,A,2 */
                    {8'hb9,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHL,A,3 */
                    {8'hc9,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHL,A,4 */
                    {8'hd9,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHL,A,5 */
                    {8'he9,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHL,A,6 */
                    {8'hf9,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SHL,A,7 */
                    {8'h88,2'bxx} : dec_alu_bitsh_adrstage = 5'h4;  /* SHL,B,0 */
                    {8'h98,2'bxx} : dec_alu_bitsh_adrstage = 5'h4;  /* SHL,B,1 */
                    {8'ha8,2'bxx} : dec_alu_bitsh_adrstage = 5'h4;  /* SHL,B,2 */
                    {8'hb8,2'bxx} : dec_alu_bitsh_adrstage = 5'h4;  /* SHL,B,3 */
                    {8'hc8,2'bxx} : dec_alu_bitsh_adrstage = 5'h4;  /* SHL,B,4 */
                    {8'hd8,2'bxx} : dec_alu_bitsh_adrstage = 5'h4;  /* SHL,B,5 */
                    {8'he8,2'bxx} : dec_alu_bitsh_adrstage = 5'h4;  /* SHL,B,6 */
                    {8'hf8,2'bxx} : dec_alu_bitsh_adrstage = 5'h4;  /* SHL,B,7 */
                    {8'h87,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHL,C,0 */
                    {8'h97,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHL,C,1 */
                    {8'ha7,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHL,C,2 */
                    {8'hb7,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHL,C,3 */
                    {8'hc7,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHL,C,4 */
                    {8'hd7,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHL,C,5 */
                    {8'he7,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHL,C,6 */
                    {8'hf7,2'bxx} : dec_alu_bitsh_adrstage = 5'h5;  /* SHL,C,7 */
                    {8'h8b,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SAR,A,0 */
                    {8'h9b,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SAR,A,1 */
                    {8'hab,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SAR,A,2 */
                    {8'hbb,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SAR,A,3 */
                    {8'hcb,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SAR,A,4 */
                    {8'hdb,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SAR,A,5 */
                    {8'heb,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SAR,A,6 */
                    {8'hfb,2'bxx} : dec_alu_bitsh_adrstage = 5'h2;  /* SAR,A,7 */
                    default : dec_alu_bitsh_adrstage = 5'h0;
                endcase
            end else begin
                    dec_alu_bitsh_adrstage = 5'h0;
            end
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_alu_bitsh <= 5'h0;
        else if(cpuen) dec_alu_bitsh <= dec_alu_bitsh_adrstage;
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*����BITEN���ѤΥǥ�������������						*/
/*------------------------------------------------------------------------------*/

    output dec_alu_biten ;
    reg    dec_alu_biten ,dec_alu_biten_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1) begin
            dec_alu_biten_adrstage = 1'b0;
        end else if(ivack == 1'b1) begin
            dec_alu_biten_adrstage = 1'b0;
        end else if(skpack == 1'b1) begin
            dec_alu_biten_adrstage = 1'b0;
        end else begin
            if(ID_stage0 == 8'h71) begin			/* MOV1, AND1, OR1, XOR1, SET1, CLR1, NOT1 */
                casex ({ID_stage1,stage_adr})  
                    {8'h01,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,saddr.0,CY */
                    {8'h11,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,saddr.1,CY */
                    {8'h21,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,saddr.2,CY */
                    {8'h31,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,saddr.3,CY */
                    {8'h41,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,saddr.4,CY */
                    {8'h51,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,saddr.5,CY */
                    {8'h61,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,saddr.6,CY */
                    {8'h71,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,saddr.7,CY */
                    {8'h09,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,sfr.0,CY */
                    {8'h19,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,sfr.1,CY */
                    {8'h29,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,sfr.2,CY */
                    {8'h39,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,sfr.3,CY */
                    {8'h49,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,sfr.4,CY */
                    {8'h59,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,sfr.5,CY */
                    {8'h69,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,sfr.6,CY */
                    {8'h79,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,sfr.7,CY */
                    {8'h81,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,[HL].0,CY */
                    {8'h91,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,[HL].1,CY */
                    {8'ha1,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,[HL].2,CY */
                    {8'hb1,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,[HL].3,CY */
                    {8'hc1,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,[HL].4,CY */
                    {8'hd1,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,[HL].5,CY */
                    {8'he1,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,[HL].6,CY */
                    {8'hf1,2'bx1} : dec_alu_biten_adrstage = 1'b1;   /* MOV1,[HL].7,CY */
                    {8'h02,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,saddr.0 */
                    {8'h12,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,saddr.1 */
                    {8'h22,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,saddr.2 */
                    {8'h32,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,saddr.3 */
                    {8'h42,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,saddr.4 */
                    {8'h52,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,saddr.5 */
                    {8'h62,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,saddr.6 */
                    {8'h72,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,saddr.7 */
                    {8'h0a,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,sfr.0 */
                    {8'h1a,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,sfr.1 */
                    {8'h2a,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,sfr.2 */
                    {8'h3a,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,sfr.3 */
                    {8'h4a,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,sfr.4 */
                    {8'h5a,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,sfr.5 */
                    {8'h6a,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,sfr.6 */
                    {8'h7a,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,sfr.7 */
                    {8'h00,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,!addr16.0 */
                    {8'h10,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,!addr16.1 */
                    {8'h20,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,!addr16.2 */
                    {8'h30,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,!addr16.3 */
                    {8'h40,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,!addr16.4 */
                    {8'h50,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,!addr16.5 */
                    {8'h60,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,!addr16.6 */
                    {8'h70,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,!addr16.7 */
                    {8'h82,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,[HL].0 */
                    {8'h92,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,[HL].1 */
                    {8'ha2,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,[HL].2 */
                    {8'hb2,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,[HL].3 */
                    {8'hc2,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,[HL].4 */
                    {8'hd2,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,[HL].5 */
                    {8'he2,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,[HL].6 */
                    {8'hf2,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* SET1,,[HL].7 */
                    {8'h03,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,saddr.0 */
                    {8'h13,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,saddr.1 */
                    {8'h23,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,saddr.2 */
                    {8'h33,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,saddr.3 */
                    {8'h43,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,saddr.4 */
                    {8'h53,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,saddr.5 */
                    {8'h63,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,saddr.6 */
                    {8'h73,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,saddr.7 */
                    {8'h0b,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,sfr.0 */
                    {8'h1b,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,sfr.1 */
                    {8'h2b,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,sfr.2 */
                    {8'h3b,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,sfr.3 */
                    {8'h4b,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,sfr.4 */
                    {8'h5b,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,sfr.5 */
                    {8'h6b,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,sfr.6 */
                    {8'h7b,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,sfr.7 */
                    {8'h08,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,!addr16.0 */
                    {8'h18,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,!addr16.1 */
                    {8'h28,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,!addr16.2 */
                    {8'h38,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,!addr16.3 */
                    {8'h48,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,!addr16.4 */
                    {8'h58,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,!addr16.5 */
                    {8'h68,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,!addr16.6 */
                    {8'h78,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,!addr16.7 */
                    {8'h83,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,[HL].0 */
                    {8'h93,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,[HL].1 */
                    {8'ha3,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,[HL].2 */
                    {8'hb3,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,[HL].3 */
                    {8'hc3,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,[HL].4 */
                    {8'hd3,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,[HL].5 */
                    {8'he3,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,[HL].6 */
                    {8'hf3,2'bx1} : dec_alu_biten_adrstage = 1'b1;  /* CLR1,,[HL].7 */
                     default : dec_alu_biten_adrstage = 1'b0;
                endcase
            end else if(ID_stage0 == 8'h31) begin                      /* SHR, SHRW, SHL, SHLW, SAR, SARW, BT, BF, BTCLR */
                casex ({ID_stage1,stage_adr})  
                    {8'h00,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,saddr.0,$addr8 */
                    {8'h10,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,saddr.1,$addr8 */
                    {8'h20,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,saddr.2,$addr8 */
                    {8'h30,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,saddr.3,$addr8 */
                    {8'h40,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,saddr.4,$addr8 */
                    {8'h50,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,saddr.5,$addr8 */
                    {8'h60,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,saddr.6,$addr8 */
                    {8'h70,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,saddr.7,$addr8 */
                    {8'h80,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,sfr.0,$addr8 */
                    {8'h90,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,sfr.1,$addr8 */
                    {8'ha0,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,sfr.2,$addr8 */
                    {8'hb0,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,sfr.3,$addr8 */
                    {8'hc0,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,sfr.4,$addr8 */
                    {8'hd0,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,sfr.5,$addr8 */
                    {8'he0,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,sfr.6,$addr8 */
                    {8'hf0,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,sfr.7,$addr8 */
                    {8'h81,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,[HL].0,$addr8 */
                    {8'h91,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,[HL].1,$addr8 */
                    {8'ha1,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,[HL].2,$addr8 */
                    {8'hb1,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,[HL].3,$addr8 */
                    {8'hc1,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,[HL].4,$addr8 */
                    {8'hd1,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,[HL].5,$addr8 */
                    {8'he1,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,[HL].6,$addr8 */
                    {8'hf1,2'b10} : dec_alu_biten_adrstage = 1'b1;  /* BTCLR,[HL].7,$addr8 */
                    default : dec_alu_biten_adrstage = 1'b0;
                endcase
            end else begin
                    dec_alu_biten_adrstage = 1'b0;
            end
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_alu_biten <= 1'b0;
        else if(cpuen) dec_alu_biten <= dec_alu_biten_adrstage;
    end

    output dec_word_access;
    reg    dec_word_access, dec_word_access_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1) begin
            dec_word_access_adrstage = 1'h0;
        end else if(ivack == 1'b1) begin
            casex ({stage_adr})  
                {2'b00} : dec_word_access_adrstage = 1'b1;  /* Interrupt */
                {2'b01} : dec_word_access_adrstage = 1'b1;  /* Interrupt */
                default : dec_word_access_adrstage = 1'h0;
            endcase
        end else if(skpack == 1'b1) begin
            dec_word_access_adrstage = 1'h0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h30,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,AX,#word */
                {8'h32,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,BC,#word */
                {8'h34,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,DE,#word */
                {8'h36,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,HL,#word */
                {8'hc9,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,saddrp,#word */
                {8'hcb,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,sfrp,#word */
                {8'had,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,AX,saddrp */
                {8'hbd,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,saddrp,AX */
                {8'hae,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,AX,sfrp */
                {8'hbe,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,sfrp,AX */
                {8'h13,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,AX,BC */
                {8'h12,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,BC,AX */
                {8'h15,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,AX,DE */
                {8'h14,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,DE,AX */
                {8'h17,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,AX,HL */
                {8'h16,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,HL,AX */
                {8'haf,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,AX,!addr16 */
                {8'hbf,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,!addr16,AX */
                {8'ha9,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,AX,[DE] */
                {8'haa,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,AX,[DE+byte] */
                {8'hb9,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,[DE],AX */
                {8'hba,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,[DE+byte],AX */
                {8'hab,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,AX,[HL] */
                {8'hac,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,AX,[HL+byte] */
                {8'hbb,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,[HL],AX */
                {8'hbc,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,[HL+byte],AX */
                {8'h59,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,AX,word[B] */
                {8'h58,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,word[B],AX */
                {8'h69,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,AX,word[C] */
                {8'h68,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,word[C],AX */
                {8'h79,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,AX,word[BC] */
                {8'h78,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,word[BC],AX */
                {8'ha8,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,AX,[SP+byte] */
                {8'hb8,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,[SP+byte],AX */
                {8'hda,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,BC,saddrp */
                {8'hdb,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,BC,!addr16 */
                {8'hea,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,DE,saddrp */
                {8'heb,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,DE,!addr16 */
                {8'hfa,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,HL,saddrp */
                {8'hfb,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MOVW,HL,!addr16 */
                {8'h33,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* XCHW,AX,BC */
                {8'h35,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* XCHW,AX,DE */
                {8'h37,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* XCHW,AX,HL */
                {8'he6,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* ONEW,,AX */
                {8'he7,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* ONEW,,BC */
                {8'hf6,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* CLRW,,AX */
                {8'hf7,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* CLRW,,BC */
                {8'h04,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* ADDW,AX,#word */
                {8'h01,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* ADDW,AX,AX */
                {8'h03,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* ADDW,AX,BC */
                {8'h05,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* ADDW,AX,DE */
                {8'h07,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* ADDW,AX,HL */
                {8'h06,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* ADDW,AX,saddrp */
                {8'h02,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* ADDW,AX,!addr16 */
                {8'h61,8'h09,2'bxx} : dec_word_access_adrstage = 1'b1;  /* ADDW,AX,[HL+byte] */
                {8'h24,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SUBW,AX,#word */
                {8'h21,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SUBW,AX,AX */
                {8'h23,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SUBW,AX,BC */
                {8'h25,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SUBW,AX,DE */
                {8'h27,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SUBW,AX,HL */
                {8'h26,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SUBW,AX,saddrp */
                {8'h22,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SUBW,AX,!addr16 */
                {8'h61,8'h29,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SUBW,AX,[HL+byte] */
                {8'h44,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* CMPW,AX,#word */
                {8'h43,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* CMPW,AX,BC */
                {8'h45,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* CMPW,AX,DE */
                {8'h47,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* CMPW,AX,HL */
                {8'h46,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* CMPW,AX,saddrp */
                {8'h42,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* CMPW,AX,!addr16 */
                {8'h61,8'h49,2'bxx} : dec_word_access_adrstage = 1'b1;  /* CMPW,AX,[HL+byte] */
                {8'hd6,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* MULU,,X */
                {8'ha1,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* INCW,,AX */
                {8'ha3,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* INCW,,BC */
                {8'ha5,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* INCW,,DE */
                {8'ha7,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* INCW,,HL */
                {8'ha6,8'hxx,2'bx0} : dec_word_access_adrstage = 1'b1;  /* INCW,,saddrp */
                {8'ha6,8'hxx,2'bx1} : dec_word_access_adrstage = 1'b1;  /* INCW,,saddrp */
                {8'ha2,8'hxx,2'bx0} : dec_word_access_adrstage = 1'b1;  /* INCW,,!addr16 */
                {8'ha2,8'hxx,2'bx1} : dec_word_access_adrstage = 1'b1;  /* INCW,,!addr16 */
                {8'h61,8'h79,2'bx0} : dec_word_access_adrstage = 1'b1;  /* INCW,,[HL+byte] */
                {8'h61,8'h79,2'bx1} : dec_word_access_adrstage = 1'b1;  /* INCW,,[HL+byte] */
                {8'hb1,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* DECW,,AX */
                {8'hb3,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* DECW,,BC */
                {8'hb5,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* DECW,,DE */
                {8'hb7,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* DECW,,HL */
                {8'hb6,8'hxx,2'bx0} : dec_word_access_adrstage = 1'b1;  /* DECW,,saddrp */
                {8'hb6,8'hxx,2'bx1} : dec_word_access_adrstage = 1'b1;  /* DECW,,saddrp */
                {8'hb2,8'hxx,2'bx0} : dec_word_access_adrstage = 1'b1;  /* DECW,,!addr16 */
                {8'hb2,8'hxx,2'bx1} : dec_word_access_adrstage = 1'b1;  /* DECW,,!addr16 */
                {8'h61,8'h89,2'bx0} : dec_word_access_adrstage = 1'b1;  /* DECW,,[HL+byte] */
                {8'h61,8'h89,2'bx1} : dec_word_access_adrstage = 1'b1;  /* DECW,,[HL+byte] */
                {8'h31,8'h0e,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHRW,AX,0 */
                {8'h31,8'h1e,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHRW,AX,1 */
                {8'h31,8'h2e,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHRW,AX,2 */
                {8'h31,8'h3e,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHRW,AX,3 */
                {8'h31,8'h4e,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHRW,AX,4 */
                {8'h31,8'h5e,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHRW,AX,5 */
                {8'h31,8'h6e,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHRW,AX,6 */
                {8'h31,8'h7e,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHRW,AX,7 */
                {8'h31,8'h8e,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHRW,AX,8 */
                {8'h31,8'h9e,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHRW,AX,9 */
                {8'h31,8'hae,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHRW,AX,10 */
                {8'h31,8'hbe,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHRW,AX,11 */
                {8'h31,8'hce,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHRW,AX,12 */
                {8'h31,8'hde,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHRW,AX,13 */
                {8'h31,8'hee,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHRW,AX,14 */
                {8'h31,8'hfe,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHRW,AX,15 */
                {8'h31,8'h0d,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,AX,0 */
                {8'h31,8'h1d,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,AX,1 */
                {8'h31,8'h2d,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,AX,2 */
                {8'h31,8'h3d,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,AX,3 */
                {8'h31,8'h4d,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,AX,4 */
                {8'h31,8'h5d,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,AX,5 */
                {8'h31,8'h6d,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,AX,6 */
                {8'h31,8'h7d,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,AX,7 */
                {8'h31,8'h8d,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,AX,8 */
                {8'h31,8'h9d,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,AX,9 */
                {8'h31,8'had,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,AX,10 */
                {8'h31,8'hbd,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,AX,11 */
                {8'h31,8'hcd,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,AX,12 */
                {8'h31,8'hdd,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,AX,13 */
                {8'h31,8'hed,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,AX,14 */
                {8'h31,8'hfd,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,AX,15 */
                {8'h31,8'h0c,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,BC,0 */
                {8'h31,8'h1c,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,BC,1 */
                {8'h31,8'h2c,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,BC,2 */
                {8'h31,8'h3c,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,BC,3 */
                {8'h31,8'h4c,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,BC,4 */
                {8'h31,8'h5c,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,BC,5 */
                {8'h31,8'h6c,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,BC,6 */
                {8'h31,8'h7c,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,BC,7 */
                {8'h31,8'h8c,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,BC,8 */
                {8'h31,8'h9c,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,BC,9 */
                {8'h31,8'hac,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,BC,10 */
                {8'h31,8'hbc,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,BC,11 */
                {8'h31,8'hcc,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,BC,12 */
                {8'h31,8'hdc,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,BC,13 */
                {8'h31,8'hec,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,BC,14 */
                {8'h31,8'hfc,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SHLW,BC,15 */
                {8'h31,8'h0f,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SARW,AX,0 */
                {8'h31,8'h1f,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SARW,AX,1 */
                {8'h31,8'h2f,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SARW,AX,2 */
                {8'h31,8'h3f,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SARW,AX,3 */
                {8'h31,8'h4f,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SARW,AX,4 */
                {8'h31,8'h5f,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SARW,AX,5 */
                {8'h31,8'h6f,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SARW,AX,6 */
                {8'h31,8'h7f,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SARW,AX,7 */
                {8'h31,8'h8f,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SARW,AX,8 */
                {8'h31,8'h9f,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SARW,AX,9 */
                {8'h31,8'haf,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SARW,AX,10 */
                {8'h31,8'hbf,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SARW,AX,11 */
                {8'h31,8'hcf,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SARW,AX,12 */
                {8'h31,8'hdf,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SARW,AX,13 */
                {8'h31,8'hef,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SARW,AX,14 */
                {8'h31,8'hff,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SARW,AX,15 */
                {8'h61,8'hee,2'bxx} : dec_word_access_adrstage = 1'b1;  /* ROLWC,AX,1 */
                {8'h61,8'hfe,2'bxx} : dec_word_access_adrstage = 1'b1;  /* ROLWC,BC,1 */
                {8'h61,8'hca,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALL,,AX */
                {8'h61,8'hda,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALL,,BC */
                {8'h61,8'hea,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALL,,DE */
                {8'h61,8'hfa,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALL,,HL */
                {8'hfe,8'hxx,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALL,,$!addr16 */
                {8'hfd,8'hxx,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALL,,!addr16 */
                {8'hfc,8'hxx,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALL,,!!addr20 */
                {8'h61,8'h84,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[0080h] */
                {8'h61,8'h94,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[0082h] */
                {8'h61,8'ha4,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[0084h] */
                {8'h61,8'hb4,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[0086h] */
                {8'h61,8'hc4,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[0088h] */
                {8'h61,8'hd4,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[008Ah] */
                {8'h61,8'he4,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[008Ch] */
                {8'h61,8'hf4,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[008Eh] */
                {8'h61,8'h85,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[0090h] */
                {8'h61,8'h95,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[0092h] */
                {8'h61,8'ha5,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[0094h] */
                {8'h61,8'hb5,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[0096h] */
                {8'h61,8'hc5,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[0098h] */
                {8'h61,8'hd5,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[009Ah] */
                {8'h61,8'he5,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[009Ch] */
                {8'h61,8'hf5,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[009Eh] */
                {8'h61,8'h86,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[00A0h] */
                {8'h61,8'h96,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[00A2h] */
                {8'h61,8'ha6,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[00A4h] */
                {8'h61,8'hb6,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[00A6h] */
                {8'h61,8'hc6,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[00A8h] */
                {8'h61,8'hd6,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[00AAh] */
                {8'h61,8'he6,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[00ACh] */
                {8'h61,8'hf6,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[00AEh] */
                {8'h61,8'h87,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[00B0h] */
                {8'h61,8'h97,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[00B2h] */
                {8'h61,8'ha7,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[00B4h] */
                {8'h61,8'hb7,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[00B6h] */
                {8'h61,8'hc7,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[00B8h] */
                {8'h61,8'hd7,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[00BAh] */
                {8'h61,8'he7,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[00BCh] */
                {8'h61,8'hf7,2'bx1} : dec_word_access_adrstage = 1'b1;  /* CALLT,,[00BEh] */
                {8'h61,8'hcc,2'bx0} : dec_word_access_adrstage = 1'b1;  /* BRK,, */
                {8'h61,8'hcc,2'bx1} : dec_word_access_adrstage = 1'b1;  /* BRK,, */
                {8'hd7,8'hxx,2'b00} : dec_word_access_adrstage = 1'b1;  /* RET,, */
                {8'h61,8'hec,2'b00} : dec_word_access_adrstage = 1'b1;  /* RETB,, */
                {8'h61,8'hec,2'b01} : dec_word_access_adrstage = 1'b1;  /* RETB,, */
                {8'h61,8'hfc,2'b00} : dec_word_access_adrstage = 1'b1;  /* RETI,, */
                {8'h61,8'hfc,2'b01} : dec_word_access_adrstage = 1'b1;  /* RETI,, */
                {8'h61,8'hdd,2'bxx} : dec_word_access_adrstage = 1'b1;  /* PUSH,,PSW */
                {8'hc1,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* PUSH,,AX */
                {8'hc3,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* PUSH,,BC */
                {8'hc5,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* PUSH,,DE */
                {8'hc7,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* PUSH,,HL */
                {8'h61,8'hcd,2'bxx} : dec_word_access_adrstage = 1'b1;  /* POP,,PSW */
                {8'hc0,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* POP,,AX */
                {8'hc2,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* POP,,BC */
                {8'hc4,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* POP,,DE */
                {8'hc6,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* POP,,HL */
                {8'h10,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* ADDW,SP,#byte */
                {8'h20,8'hxx,2'bxx} : dec_word_access_adrstage = 1'b1;  /* SUBW,SP,#byte */
                {8'hff,8'hxx,2'bx0} : dec_word_access_adrstage = 1'b1;  /* SOFT,,BREAK */
                {8'hff,8'hxx,2'bx1} : dec_word_access_adrstage = 1'b1;  /* SOFT,,BREAK */
                {8'h61,8'ha1,2'bx0} : dec_word_access_adrstage = 1'b1;  /* SOFT2,,BREAK */
                {8'h61,8'ha1,2'bx1} : dec_word_access_adrstage = 1'b1;  /* SOFT2,,BREAK */
                {8'h61,8'hb1,2'bx0} : dec_word_access_adrstage = 1'b1;  /* SOFT3,,BREAK */
                {8'h61,8'hb1,2'bx1} : dec_word_access_adrstage = 1'b1;  /* SOFT3,,BREAK */
                {8'h61,8'hc1,2'bx0} : dec_word_access_adrstage = 1'b1;  /* SOFT4,,BREAK */
                {8'h61,8'hc1,2'bx1} : dec_word_access_adrstage = 1'b1;  /* SOFT4,,BREAK */
                default : dec_word_access_adrstage = 1'h0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_word_access <= 1'b0;
        else if(cpuen) dec_word_access <= dec_word_access_adrstage;
    end
    output dec_xch_byte;
    reg    dec_xch_byte, dec_xch_byte_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_xch_byte_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h08,8'hxx,2'bxx} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,X */
                {8'h61,8'h8a,2'bxx} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,C */
                {8'h61,8'h8b,2'bxx} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,B */
                {8'h61,8'h8c,2'bxx} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,E */
                {8'h61,8'h8d,2'bxx} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,D */
                {8'h61,8'h8e,2'bxx} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,L */
                {8'h61,8'h8f,2'bxx} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,H */
                {8'h61,8'ha8,2'bx1} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,saddr */
                {8'h61,8'hab,2'bx1} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,sfr */
                {8'h61,8'haa,2'bx1} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,!addr16 */
                {8'h61,8'hae,2'bx1} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,[DE] */
                {8'h61,8'haf,2'bx1} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,[DE+byte] */
                {8'h61,8'hac,2'bx1} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,[HL] */
                {8'h61,8'had,2'bx1} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,[HL+byte] */
                {8'h61,8'hb9,2'bx1} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,[HL+B] */
                {8'h61,8'ha9,2'bx1} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,[HL+C] */
                {8'h61,8'h88,2'bxx} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,X */
                {8'h61,8'h98,2'bxx} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,X */
                {8'h61,8'h99,2'bxx} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,X */
                {8'h61,8'h9a,2'bxx} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,C */
                {8'h61,8'h9b,2'bxx} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,B */
                {8'h61,8'h9c,2'bxx} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,E */
                {8'h61,8'h9d,2'bxx} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,D */
                {8'h61,8'h9e,2'bxx} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,L */
                {8'h61,8'h9f,2'bxx} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,H */
                {8'h61,8'hbb,2'bx1} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,sfr */
                {8'h61,8'hba,2'bx1} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,!addr16 */
                {8'h61,8'hbe,2'bx1} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,[DE] */
                {8'h61,8'hbf,2'bx1} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,[DE+byte] */
                {8'h61,8'hbc,2'bx1} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,[HL] */
                {8'h61,8'hbd,2'bx1} : dec_xch_byte_adrstage = 1'b1;  /* XCH,A,[HL+byte] */
                default : dec_xch_byte_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_xch_byte <= 1'b0;
        else if(cpuen) dec_xch_byte <= dec_xch_byte_adrstage;
    end
    output dec_xchw_bc;
    reg    dec_xchw_bc, dec_xchw_bc_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_xchw_bc_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h33,8'hxx,2'bxx} : dec_xchw_bc_adrstage = 1'b1;  /* XCHW,AX,BC */
                default : dec_xchw_bc_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_xchw_bc <= 1'b0;
        else if(cpuen) dec_xchw_bc <= dec_xchw_bc_adrstage;
    end
    output dec_xchw_de;
    reg    dec_xchw_de, dec_xchw_de_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_xchw_de_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h35,8'hxx,2'bxx} : dec_xchw_de_adrstage = 1'b1;  /* XCHW,AX,DE */
                default : dec_xchw_de_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_xchw_de <= 1'b0;
        else if(cpuen) dec_xchw_de <= dec_xchw_de_adrstage;
    end
    output dec_xchw_hl;
    reg    dec_xchw_hl, dec_xchw_hl_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_xchw_hl_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h37,8'hxx,2'bxx} : dec_xchw_hl_adrstage = 1'b1;  /* XCHW,AX,HL */
                default : dec_xchw_hl_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_xchw_hl <= 1'b0;
        else if(cpuen) dec_xchw_hl <= dec_xchw_hl_adrstage;
    end
    output dec_SP_enable;
    reg    dec_SP_enable, dec_SP_enable_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1|| skpack == 1'b1) begin
            dec_SP_enable_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h10,8'hxx,2'bxx} : dec_SP_enable_adrstage = 1'b1;  /* ADDW,SP,#byte */
                {8'h20,8'hxx,2'bxx} : dec_SP_enable_adrstage = 1'b1;  /* SUBW,SP,#byte */
                default : dec_SP_enable_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_SP_enable <= 1'b0;
        else if(cpuen) dec_SP_enable <= dec_SP_enable_adrstage;
    end
    output dec_A_enable;
    reg    dec_A_enable, dec_A_enable_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1|| skpack == 1'b1) begin
            dec_A_enable_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h51,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV,A,#byte */
                {8'h60,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV,A,X */
                {8'h62,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV,A,C */
                {8'h63,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV,A,B */
                {8'h64,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV,A,E */
                {8'h65,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV,A,D */
                {8'h66,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV,A,L */
                {8'h67,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV,A,H */
                {8'h8d,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV,A,saddr */
                {8'h8e,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV,A,sfr */
                {8'h8f,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV,A,!addr16 */
                {8'h89,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV,A,[DE] */
                {8'h8a,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV,A,[DE+byte] */
                {8'h8b,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV,A,[HL] */
                {8'h8c,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV,A,[HL+byte] */
                {8'h61,8'hc9,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV,A,[HL+B] */
                {8'h61,8'he9,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV,A,[HL+C] */
                {8'h09,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV,A,word[B] */
                {8'h29,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV,A,word[C] */
                {8'h49,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV,A,word[BC] */
                {8'h88,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV,A,[SP+byte] */
                {8'h08,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,X */
                {8'h61,8'h8a,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,C */
                {8'h61,8'h8b,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,B */
                {8'h61,8'h8c,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,E */
                {8'h61,8'h8d,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,D */
                {8'h61,8'h8e,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,L */
                {8'h61,8'h8f,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,H */
                {8'h61,8'ha8,2'bx1} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,saddr */
                {8'h61,8'hab,2'bx1} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,sfr */
                {8'h61,8'haa,2'bx1} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,!addr16 */
                {8'h61,8'hae,2'bx1} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,[DE] */
                {8'h61,8'haf,2'bx1} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,[DE+byte] */
                {8'h61,8'hac,2'bx1} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,[HL] */
                {8'h61,8'had,2'bx1} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,[HL+byte] */
                {8'h61,8'hb9,2'bx1} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,[HL+B] */
                {8'h61,8'ha9,2'bx1} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,[HL+C] */
                {8'he1,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ONEB,,A */
                {8'hf1,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* CLRB,,A */
                {8'h30,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOVW,AX,#word */
                {8'had,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOVW,AX,saddrp */
                {8'hae,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOVW,AX,sfrp */
                {8'h13,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOVW,AX,BC */
                {8'h15,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOVW,AX,DE */
                {8'h17,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOVW,AX,HL */
                {8'haf,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOVW,AX,!addr16 */
                {8'ha9,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOVW,AX,[DE] */
                {8'haa,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOVW,AX,[DE+byte] */
                {8'hab,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOVW,AX,[HL] */
                {8'hac,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOVW,AX,[HL+byte] */
                {8'h59,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOVW,AX,word[B] */
                {8'h69,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOVW,AX,word[C] */
                {8'h79,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOVW,AX,word[BC] */
                {8'ha8,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOVW,AX,[SP+byte] */
                {8'h33,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XCHW,AX,BC */
                {8'h35,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XCHW,AX,DE */
                {8'h37,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XCHW,AX,HL */
                {8'he6,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ONEW,,AX */
                {8'hf6,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* CLRW,,AX */
                {8'h0c,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADD,A,#byte */
                {8'h61,8'h08,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADD,A,X */
                {8'h61,8'h0a,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADD,A,C */
                {8'h61,8'h0b,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADD,A,B */
                {8'h61,8'h0c,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADD,A,E */
                {8'h61,8'h0d,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADD,A,D */
                {8'h61,8'h0e,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADD,A,L */
                {8'h61,8'h0f,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADD,A,H */
                {8'h61,8'h01,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADD,A,A */
                {8'h0b,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADD,A,saddr */
                {8'h0f,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADD,A,!addr16 */
                {8'h0d,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADD,A,[HL] */
                {8'h0e,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADD,A,[HL+byte] */
                {8'h61,8'h80,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADD,A,[HL+B] */
                {8'h61,8'h82,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADD,A,[HL+C] */
                {8'h1c,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDC,A,#byte */
                {8'h61,8'h18,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDC,A,X */
                {8'h61,8'h1a,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDC,A,C */
                {8'h61,8'h1b,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDC,A,B */
                {8'h61,8'h1c,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDC,A,E */
                {8'h61,8'h1d,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDC,A,D */
                {8'h61,8'h1e,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDC,A,L */
                {8'h61,8'h1f,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDC,A,H */
                {8'h61,8'h11,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDC,A,A */
                {8'h1b,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDC,A,saddr */
                {8'h1f,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDC,A,!addr16 */
                {8'h1d,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDC,A,[HL] */
                {8'h1e,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDC,A,[HL+byte] */
                {8'h61,8'h90,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDC,A,[HL+B] */
                {8'h61,8'h92,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDC,A,[HL+C] */
                {8'h2c,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUB,A,#byte */
                {8'h61,8'h28,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUB,A,X */
                {8'h61,8'h2a,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUB,A,C */
                {8'h61,8'h2b,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUB,A,B */
                {8'h61,8'h2c,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUB,A,E */
                {8'h61,8'h2d,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUB,A,D */
                {8'h61,8'h2e,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUB,A,L */
                {8'h61,8'h2f,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUB,A,H */
                {8'h61,8'h21,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUB,A,A */
                {8'h2b,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUB,A,saddr */
                {8'h2f,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUB,A,!addr16 */
                {8'h2d,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUB,A,[HL] */
                {8'h2e,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUB,A,[HL+byte] */
                {8'h61,8'ha0,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUB,A,[HL+B] */
                {8'h61,8'ha2,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUB,A,[HL+C] */
                {8'h3c,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBC,A,#byte */
                {8'h61,8'h38,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBC,A,X */
                {8'h61,8'h3a,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBC,A,C */
                {8'h61,8'h3b,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBC,A,B */
                {8'h61,8'h3c,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBC,A,E */
                {8'h61,8'h3d,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBC,A,D */
                {8'h61,8'h3e,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBC,A,L */
                {8'h61,8'h3f,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBC,A,H */
                {8'h61,8'h31,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBC,A,A */
                {8'h3b,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBC,A,saddr */
                {8'h3f,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBC,A,!addr16 */
                {8'h3d,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBC,A,[HL] */
                {8'h3e,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBC,A,[HL+byte] */
                {8'h61,8'hb0,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBC,A,[HL+B] */
                {8'h61,8'hb2,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBC,A,[HL+C] */
                {8'h5c,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* AND,A,#byte */
                {8'h61,8'h58,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* AND,A,X */
                {8'h61,8'h5a,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* AND,A,C */
                {8'h61,8'h5b,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* AND,A,B */
                {8'h61,8'h5c,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* AND,A,E */
                {8'h61,8'h5d,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* AND,A,D */
                {8'h61,8'h5e,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* AND,A,L */
                {8'h61,8'h5f,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* AND,A,H */
                {8'h61,8'h51,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* AND,A,A */
                {8'h5b,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* AND,A,saddr */
                {8'h5f,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* AND,A,!addr16 */
                {8'h5d,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* AND,A,[HL] */
                {8'h5e,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* AND,A,[HL+byte] */
                {8'h61,8'hd0,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* AND,A,[HL+B] */
                {8'h61,8'hd2,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* AND,A,[HL+C] */
                {8'h6c,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* OR,A,#byte */
                {8'h61,8'h68,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* OR,A,X */
                {8'h61,8'h6a,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* OR,A,C */
                {8'h61,8'h6b,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* OR,A,B */
                {8'h61,8'h6c,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* OR,A,E */
                {8'h61,8'h6d,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* OR,A,D */
                {8'h61,8'h6e,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* OR,A,L */
                {8'h61,8'h6f,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* OR,A,H */
                {8'h61,8'h61,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* OR,A,A */
                {8'h6b,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* OR,A,saddr */
                {8'h6f,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* OR,A,!addr16 */
                {8'h6d,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* OR,A,[HL] */
                {8'h6e,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* OR,A,[HL+byte] */
                {8'h61,8'he0,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* OR,A,[HL+B] */
                {8'h61,8'he2,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* OR,A,[HL+C] */
                {8'h7c,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XOR,A,#byte */
                {8'h61,8'h78,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XOR,A,X */
                {8'h61,8'h7a,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XOR,A,C */
                {8'h61,8'h7b,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XOR,A,B */
                {8'h61,8'h7c,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XOR,A,E */
                {8'h61,8'h7d,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XOR,A,D */
                {8'h61,8'h7e,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XOR,A,L */
                {8'h61,8'h7f,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XOR,A,H */
                {8'h61,8'h71,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XOR,A,A */
                {8'h7b,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XOR,A,saddr */
                {8'h7f,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XOR,A,!addr16 */
                {8'h7d,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XOR,A,[HL] */
                {8'h7e,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XOR,A,[HL+byte] */
                {8'h61,8'hf0,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XOR,A,[HL+B] */
                {8'h61,8'hf2,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XOR,A,[HL+C] */
                {8'h04,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDW,AX,#word */
                {8'h01,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDW,AX,AX */
                {8'h03,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDW,AX,BC */
                {8'h05,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDW,AX,DE */
                {8'h07,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDW,AX,HL */
                {8'h06,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDW,AX,saddrp */
                {8'h02,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDW,AX,!addr16 */
                {8'h61,8'h09,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDW,AX,[HL+byte] */
                {8'h24,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBW,AX,#word */
                {8'h21,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBW,AX,AX */
                {8'h23,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBW,AX,BC */
                {8'h25,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBW,AX,DE */
                {8'h27,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBW,AX,HL */
                {8'h26,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBW,AX,saddrp */
                {8'h22,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBW,AX,!addr16 */
                {8'h61,8'h29,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBW,AX,[HL+byte] */
                {8'hd6,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MULU,,X */
                {8'h81,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* INC,,A */
                {8'h91,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* DEC,,A */
                {8'ha1,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* INCW,,AX */
                {8'hb1,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* DECW,,AX */
                {8'h31,8'h0a,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHR,A,0 */
                {8'h31,8'h1a,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHR,A,1 */
                {8'h31,8'h2a,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHR,A,2 */
                {8'h31,8'h3a,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHR,A,3 */
                {8'h31,8'h4a,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHR,A,4 */
                {8'h31,8'h5a,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHR,A,5 */
                {8'h31,8'h6a,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHR,A,6 */
                {8'h31,8'h7a,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHR,A,7 */
                {8'h31,8'h0e,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHRW,AX,0 */
                {8'h31,8'h1e,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHRW,AX,1 */
                {8'h31,8'h2e,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHRW,AX,2 */
                {8'h31,8'h3e,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHRW,AX,3 */
                {8'h31,8'h4e,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHRW,AX,4 */
                {8'h31,8'h5e,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHRW,AX,5 */
                {8'h31,8'h6e,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHRW,AX,6 */
                {8'h31,8'h7e,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHRW,AX,7 */
                {8'h31,8'h8e,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHRW,AX,8 */
                {8'h31,8'h9e,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHRW,AX,9 */
                {8'h31,8'hae,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHRW,AX,10 */
                {8'h31,8'hbe,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHRW,AX,11 */
                {8'h31,8'hce,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHRW,AX,12 */
                {8'h31,8'hde,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHRW,AX,13 */
                {8'h31,8'hee,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHRW,AX,14 */
                {8'h31,8'hfe,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHRW,AX,15 */
                {8'h31,8'h09,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHL,A,0 */
                {8'h31,8'h19,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHL,A,1 */
                {8'h31,8'h29,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHL,A,2 */
                {8'h31,8'h39,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHL,A,3 */
                {8'h31,8'h49,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHL,A,4 */
                {8'h31,8'h59,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHL,A,5 */
                {8'h31,8'h69,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHL,A,6 */
                {8'h31,8'h79,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHL,A,7 */
                {8'h31,8'h0d,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHLW,AX,0 */
                {8'h31,8'h1d,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHLW,AX,1 */
                {8'h31,8'h2d,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHLW,AX,2 */
                {8'h31,8'h3d,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHLW,AX,3 */
                {8'h31,8'h4d,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHLW,AX,4 */
                {8'h31,8'h5d,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHLW,AX,5 */
                {8'h31,8'h6d,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHLW,AX,6 */
                {8'h31,8'h7d,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHLW,AX,7 */
                {8'h31,8'h8d,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHLW,AX,8 */
                {8'h31,8'h9d,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHLW,AX,9 */
                {8'h31,8'had,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHLW,AX,10 */
                {8'h31,8'hbd,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHLW,AX,11 */
                {8'h31,8'hcd,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHLW,AX,12 */
                {8'h31,8'hdd,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHLW,AX,13 */
                {8'h31,8'hed,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHLW,AX,14 */
                {8'h31,8'hfd,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHLW,AX,15 */
                {8'h31,8'h0b,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SAR,A,0 */
                {8'h31,8'h1b,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SAR,A,1 */
                {8'h31,8'h2b,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SAR,A,2 */
                {8'h31,8'h3b,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SAR,A,3 */
                {8'h31,8'h4b,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SAR,A,4 */
                {8'h31,8'h5b,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SAR,A,5 */
                {8'h31,8'h6b,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SAR,A,6 */
                {8'h31,8'h7b,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SAR,A,7 */
                {8'h31,8'h0f,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SARW,AX,0 */
                {8'h31,8'h1f,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SARW,AX,1 */
                {8'h31,8'h2f,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SARW,AX,2 */
                {8'h31,8'h3f,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SARW,AX,3 */
                {8'h31,8'h4f,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SARW,AX,4 */
                {8'h31,8'h5f,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SARW,AX,5 */
                {8'h31,8'h6f,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SARW,AX,6 */
                {8'h31,8'h7f,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SARW,AX,7 */
                {8'h31,8'h8f,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SARW,AX,8 */
                {8'h31,8'h9f,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SARW,AX,9 */
                {8'h31,8'haf,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SARW,AX,10 */
                {8'h31,8'hbf,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SARW,AX,11 */
                {8'h31,8'hcf,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SARW,AX,12 */
                {8'h31,8'hdf,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SARW,AX,13 */
                {8'h31,8'hef,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SARW,AX,14 */
                {8'h31,8'hff,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SARW,AX,15 */
                {8'h61,8'hdb,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ROR,A,1 */
                {8'h61,8'heb,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ROL,A,1 */
                {8'h61,8'hfb,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* RORC,A,1 */
                {8'h61,8'hdc,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ROLC,A,1 */
                {8'h61,8'hee,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ROLWC,AX,1 */
                {8'h71,8'h89,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV1,A.0,CY */
                {8'h71,8'h99,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV1,A.1,CY */
                {8'h71,8'ha9,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV1,A.2,CY */
                {8'h71,8'hb9,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV1,A.3,CY */
                {8'h71,8'hc9,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV1,A.4,CY */
                {8'h71,8'hd9,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV1,A.5,CY */
                {8'h71,8'he9,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV1,A.6,CY */
                {8'h71,8'hf9,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* MOV1,A.7,CY */
                {8'h71,8'h8a,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SET1,,A.0 */
                {8'h71,8'h9a,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SET1,,A.1 */
                {8'h71,8'haa,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SET1,,A.2 */
                {8'h71,8'hba,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SET1,,A.3 */
                {8'h71,8'hca,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SET1,,A.4 */
                {8'h71,8'hda,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SET1,,A.5 */
                {8'h71,8'hea,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SET1,,A.6 */
                {8'h71,8'hfa,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SET1,,A.7 */
                {8'h71,8'h8b,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* CLR1,,A.0 */
                {8'h71,8'h9b,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* CLR1,,A.1 */
                {8'h71,8'hab,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* CLR1,,A.2 */
                {8'h71,8'hbb,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* CLR1,,A.3 */
                {8'h71,8'hcb,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* CLR1,,A.4 */
                {8'h71,8'hdb,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* CLR1,,A.5 */
                {8'h71,8'heb,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* CLR1,,A.6 */
                {8'h71,8'hfb,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* CLR1,,A.7 */
                {8'hc0,8'hxx,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* POP,,AX */
                {8'h31,8'h01,2'b10} : dec_A_enable_adrstage = 1'b1;  /* BTCLR,A.0,$addr8 */
                {8'h31,8'h11,2'b10} : dec_A_enable_adrstage = 1'b1;  /* BTCLR,A.1,$addr8 */
                {8'h31,8'h21,2'b10} : dec_A_enable_adrstage = 1'b1;  /* BTCLR,A.2,$addr8 */
                {8'h31,8'h31,2'b10} : dec_A_enable_adrstage = 1'b1;  /* BTCLR,A.3,$addr8 */
                {8'h31,8'h41,2'b10} : dec_A_enable_adrstage = 1'b1;  /* BTCLR,A.4,$addr8 */
                {8'h31,8'h51,2'b10} : dec_A_enable_adrstage = 1'b1;  /* BTCLR,A.5,$addr8 */
                {8'h31,8'h61,2'b10} : dec_A_enable_adrstage = 1'b1;  /* BTCLR,A.6,$addr8 */
                {8'h31,8'h71,2'b10} : dec_A_enable_adrstage = 1'b1;  /* BTCLR,A.7,$addr8 */
                {8'h61,8'h88,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,X */
                {8'h61,8'h98,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,X */
                {8'h61,8'h99,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,X */
                {8'h61,8'h9a,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,C */
                {8'h61,8'h9b,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,B */
                {8'h61,8'h9c,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,E */
                {8'h61,8'h9d,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,D */
                {8'h61,8'h9e,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,L */
                {8'h61,8'h9f,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,H */
                {8'h61,8'hbb,2'bx1} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,sfr */
                {8'h61,8'hba,2'bx1} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,!addr16 */
                {8'h61,8'hbe,2'bx1} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,[DE] */
                {8'h61,8'hbf,2'bx1} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,[DE+byte] */
                {8'h61,8'hbc,2'bx1} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,[HL] */
                {8'h61,8'hbd,2'bx1} : dec_A_enable_adrstage = 1'b1;  /* XCH,A,[HL+byte] */
                {8'h61,8'h19,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDC,A,A */
                {8'h61,8'h39,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBC,A,A */
                {8'h61,8'hd1,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* AND,A,[HL+B] */
                {8'h61,8'he1,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* OR,A,[HL+B] */
                {8'h61,8'hf1,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* XOR,A,[HL+B] */
                {8'h61,8'h83,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADD,A,[HL+C] */
                {8'h61,8'h93,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* ADDC,A,[HL+C] */
                {8'h61,8'ha3,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUB,A,[HL+C] */
                {8'h61,8'hb3,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SUBC,A,[HL+C] */
                {8'h31,8'h8a,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHR,A,0 */
                {8'h31,8'h9a,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHR,A,1 */
                {8'h31,8'haa,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHR,A,2 */
                {8'h31,8'hba,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHR,A,3 */
                {8'h31,8'hca,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHR,A,4 */
                {8'h31,8'hda,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHR,A,5 */
                {8'h31,8'hea,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHR,A,6 */
                {8'h31,8'hfa,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHR,A,7 */
                {8'h31,8'h89,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHL,A,0 */
                {8'h31,8'h99,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHL,A,1 */
                {8'h31,8'ha9,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHL,A,2 */
                {8'h31,8'hb9,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHL,A,3 */
                {8'h31,8'hc9,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHL,A,4 */
                {8'h31,8'hd9,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHL,A,5 */
                {8'h31,8'he9,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHL,A,6 */
                {8'h31,8'hf9,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SHL,A,7 */
                {8'h31,8'h8b,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SAR,A,0 */
                {8'h31,8'h9b,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SAR,A,1 */
                {8'h31,8'hab,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SAR,A,2 */
                {8'h31,8'hbb,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SAR,A,3 */
                {8'h31,8'hcb,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SAR,A,4 */
                {8'h31,8'hdb,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SAR,A,5 */
                {8'h31,8'heb,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SAR,A,6 */
                {8'h31,8'hfb,2'bxx} : dec_A_enable_adrstage = 1'b1;  /* SAR,A,7 */
                default : dec_A_enable_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_A_enable <= 1'b0;
        else if(cpuen) dec_A_enable <= dec_A_enable_adrstage;
    end
    output dec_X_enable;
    reg    dec_X_enable, dec_X_enable_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1|| skpack == 1'b1) begin
            dec_X_enable_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h50,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* MOV,X,#byte */
                {8'h70,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* MOV,X,A */
                {8'hd8,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* MOV,X,saddr */
                {8'hd9,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* MOV,X,!addr16 */
                {8'h08,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* XCH,A,X */
                {8'he0,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* ONEB,,X */
                {8'hf0,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* CLRB,,X */
                {8'h30,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* MOVW,AX,#word */
                {8'had,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* MOVW,AX,saddrp */
                {8'hae,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* MOVW,AX,sfrp */
                {8'h13,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* MOVW,AX,BC */
                {8'h15,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* MOVW,AX,DE */
                {8'h17,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* MOVW,AX,HL */
                {8'haf,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* MOVW,AX,!addr16 */
                {8'ha9,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* MOVW,AX,[DE] */
                {8'haa,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* MOVW,AX,[DE+byte] */
                {8'hab,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* MOVW,AX,[HL] */
                {8'hac,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* MOVW,AX,[HL+byte] */
                {8'h59,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* MOVW,AX,word[B] */
                {8'h69,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* MOVW,AX,word[C] */
                {8'h79,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* MOVW,AX,word[BC] */
                {8'ha8,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* MOVW,AX,[SP+byte] */
                {8'h33,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* XCHW,AX,BC */
                {8'h35,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* XCHW,AX,DE */
                {8'h37,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* XCHW,AX,HL */
                {8'he6,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* ONEW,,AX */
                {8'hf6,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* CLRW,,AX */
                {8'h61,8'h00,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* ADD,X,A */
                {8'h61,8'h10,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* ADDC,X,A */
                {8'h61,8'h20,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SUB,X,A */
                {8'h61,8'h30,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SUBC,X,A */
                {8'h61,8'h50,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* AND,X,A */
                {8'h61,8'h60,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* OR,X,A */
                {8'h61,8'h70,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* XOR,X,A */
                {8'h04,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* ADDW,AX,#word */
                {8'h01,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* ADDW,AX,AX */
                {8'h03,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* ADDW,AX,BC */
                {8'h05,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* ADDW,AX,DE */
                {8'h07,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* ADDW,AX,HL */
                {8'h06,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* ADDW,AX,saddrp */
                {8'h02,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* ADDW,AX,!addr16 */
                {8'h61,8'h09,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* ADDW,AX,[HL+byte] */
                {8'h24,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SUBW,AX,#word */
                {8'h21,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SUBW,AX,AX */
                {8'h23,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SUBW,AX,BC */
                {8'h25,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SUBW,AX,DE */
                {8'h27,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SUBW,AX,HL */
                {8'h26,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SUBW,AX,saddrp */
                {8'h22,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SUBW,AX,!addr16 */
                {8'h61,8'h29,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SUBW,AX,[HL+byte] */
                {8'hd6,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* MULU,,X */
                {8'h80,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* INC,,X */
                {8'h90,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* DEC,,X */
                {8'ha1,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* INCW,,AX */
                {8'hb1,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* DECW,,AX */
                {8'h31,8'h0e,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHRW,AX,0 */
                {8'h31,8'h1e,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHRW,AX,1 */
                {8'h31,8'h2e,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHRW,AX,2 */
                {8'h31,8'h3e,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHRW,AX,3 */
                {8'h31,8'h4e,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHRW,AX,4 */
                {8'h31,8'h5e,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHRW,AX,5 */
                {8'h31,8'h6e,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHRW,AX,6 */
                {8'h31,8'h7e,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHRW,AX,7 */
                {8'h31,8'h8e,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHRW,AX,8 */
                {8'h31,8'h9e,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHRW,AX,9 */
                {8'h31,8'hae,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHRW,AX,10 */
                {8'h31,8'hbe,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHRW,AX,11 */
                {8'h31,8'hce,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHRW,AX,12 */
                {8'h31,8'hde,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHRW,AX,13 */
                {8'h31,8'hee,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHRW,AX,14 */
                {8'h31,8'hfe,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHRW,AX,15 */
                {8'h31,8'h0d,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHLW,AX,0 */
                {8'h31,8'h1d,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHLW,AX,1 */
                {8'h31,8'h2d,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHLW,AX,2 */
                {8'h31,8'h3d,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHLW,AX,3 */
                {8'h31,8'h4d,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHLW,AX,4 */
                {8'h31,8'h5d,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHLW,AX,5 */
                {8'h31,8'h6d,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHLW,AX,6 */
                {8'h31,8'h7d,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHLW,AX,7 */
                {8'h31,8'h8d,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHLW,AX,8 */
                {8'h31,8'h9d,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHLW,AX,9 */
                {8'h31,8'had,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHLW,AX,10 */
                {8'h31,8'hbd,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHLW,AX,11 */
                {8'h31,8'hcd,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHLW,AX,12 */
                {8'h31,8'hdd,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHLW,AX,13 */
                {8'h31,8'hed,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHLW,AX,14 */
                {8'h31,8'hfd,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SHLW,AX,15 */
                {8'h31,8'h0f,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SARW,AX,0 */
                {8'h31,8'h1f,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SARW,AX,1 */
                {8'h31,8'h2f,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SARW,AX,2 */
                {8'h31,8'h3f,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SARW,AX,3 */
                {8'h31,8'h4f,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SARW,AX,4 */
                {8'h31,8'h5f,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SARW,AX,5 */
                {8'h31,8'h6f,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SARW,AX,6 */
                {8'h31,8'h7f,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SARW,AX,7 */
                {8'h31,8'h8f,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SARW,AX,8 */
                {8'h31,8'h9f,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SARW,AX,9 */
                {8'h31,8'haf,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SARW,AX,10 */
                {8'h31,8'hbf,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SARW,AX,11 */
                {8'h31,8'hcf,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SARW,AX,12 */
                {8'h31,8'hdf,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SARW,AX,13 */
                {8'h31,8'hef,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SARW,AX,14 */
                {8'h31,8'hff,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* SARW,AX,15 */
                {8'h61,8'hee,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* ROLWC,AX,1 */
                {8'hc0,8'hxx,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* POP,,AX */
                {8'h61,8'h88,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* XCH,A,X */
                {8'h61,8'h98,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* XCH,A,X */
                {8'h61,8'h99,2'bxx} : dec_X_enable_adrstage = 1'b1;  /* XCH,A,X */
                default : dec_X_enable_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_X_enable <= 1'b0;
        else if(cpuen) dec_X_enable <= dec_X_enable_adrstage;
    end
    output dec_B_enable;
    reg    dec_B_enable, dec_B_enable_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1|| skpack == 1'b1) begin
            dec_B_enable_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h53,8'hxx,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* MOV,B,#byte */
                {8'h73,8'hxx,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* MOV,B,A */
                {8'he8,8'hxx,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* MOV,B,saddr */
                {8'he9,8'hxx,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* MOV,B,!addr16 */
                {8'h61,8'h8b,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* XCH,A,B */
                {8'he3,8'hxx,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* ONEB,,B */
                {8'hf3,8'hxx,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* CLRB,,B */
                {8'h32,8'hxx,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* MOVW,BC,#word */
                {8'h12,8'hxx,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* MOVW,BC,AX */
                {8'hda,8'hxx,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* MOVW,BC,saddrp */
                {8'hdb,8'hxx,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* MOVW,BC,!addr16 */
                {8'h33,8'hxx,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* XCHW,AX,BC */
                {8'he7,8'hxx,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* ONEW,,BC */
                {8'hf7,8'hxx,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* CLRW,,BC */
                {8'h61,8'h03,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* ADD,B,A */
                {8'h61,8'h13,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* ADDC,B,A */
                {8'h61,8'h23,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SUB,B,A */
                {8'h61,8'h33,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SUBC,B,A */
                {8'h61,8'h53,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* AND,B,A */
                {8'h61,8'h63,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* OR,B,A */
                {8'h61,8'h73,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* XOR,B,A */
                {8'h83,8'hxx,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* INC,,B */
                {8'h93,8'hxx,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* DEC,,B */
                {8'ha3,8'hxx,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* INCW,,BC */
                {8'hb3,8'hxx,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* DECW,,BC */
                {8'h31,8'h08,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHL,B,0 */
                {8'h31,8'h18,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHL,B,1 */
                {8'h31,8'h28,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHL,B,2 */
                {8'h31,8'h38,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHL,B,3 */
                {8'h31,8'h48,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHL,B,4 */
                {8'h31,8'h58,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHL,B,5 */
                {8'h31,8'h68,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHL,B,6 */
                {8'h31,8'h78,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHL,B,7 */
                {8'h31,8'h0c,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHLW,BC,0 */
                {8'h31,8'h1c,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHLW,BC,1 */
                {8'h31,8'h2c,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHLW,BC,2 */
                {8'h31,8'h3c,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHLW,BC,3 */
                {8'h31,8'h4c,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHLW,BC,4 */
                {8'h31,8'h5c,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHLW,BC,5 */
                {8'h31,8'h6c,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHLW,BC,6 */
                {8'h31,8'h7c,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHLW,BC,7 */
                {8'h31,8'h8c,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHLW,BC,8 */
                {8'h31,8'h9c,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHLW,BC,9 */
                {8'h31,8'hac,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHLW,BC,10 */
                {8'h31,8'hbc,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHLW,BC,11 */
                {8'h31,8'hcc,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHLW,BC,12 */
                {8'h31,8'hdc,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHLW,BC,13 */
                {8'h31,8'hec,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHLW,BC,14 */
                {8'h31,8'hfc,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHLW,BC,15 */
                {8'h61,8'hfe,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* ROLWC,BC,1 */
                {8'hc2,8'hxx,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* POP,,BC */
                {8'h61,8'h9b,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* XCH,A,B */
                {8'h31,8'h88,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHL,B,0 */
                {8'h31,8'h98,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHL,B,1 */
                {8'h31,8'ha8,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHL,B,2 */
                {8'h31,8'hb8,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHL,B,3 */
                {8'h31,8'hc8,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHL,B,4 */
                {8'h31,8'hd8,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHL,B,5 */
                {8'h31,8'he8,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHL,B,6 */
                {8'h31,8'hf8,2'bxx} : dec_B_enable_adrstage = 1'b1;  /* SHL,B,7 */
                default : dec_B_enable_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_B_enable <= 1'b0;
        else if(cpuen) dec_B_enable <= dec_B_enable_adrstage;
    end
    output dec_C_enable;
    reg    dec_C_enable, dec_C_enable_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1|| skpack == 1'b1) begin
            dec_C_enable_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h52,8'hxx,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* MOV,C,#byte */
                {8'h72,8'hxx,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* MOV,C,A */
                {8'hf8,8'hxx,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* MOV,C,saddr */
                {8'hf9,8'hxx,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* MOV,C,!addr16 */
                {8'h61,8'h8a,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* XCH,A,C */
                {8'he2,8'hxx,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* ONEB,,C */
                {8'hf2,8'hxx,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* CLRB,,C */
                {8'h32,8'hxx,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* MOVW,BC,#word */
                {8'h12,8'hxx,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* MOVW,BC,AX */
                {8'hda,8'hxx,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* MOVW,BC,saddrp */
                {8'hdb,8'hxx,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* MOVW,BC,!addr16 */
                {8'h33,8'hxx,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* XCHW,AX,BC */
                {8'he7,8'hxx,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* ONEW,,BC */
                {8'hf7,8'hxx,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* CLRW,,BC */
                {8'h61,8'h02,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* ADD,C,A */
                {8'h61,8'h12,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* ADDC,C,A */
                {8'h61,8'h22,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SUB,C,A */
                {8'h61,8'h32,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SUBC,C,A */
                {8'h61,8'h52,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* AND,C,A */
                {8'h61,8'h62,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* OR,C,A */
                {8'h61,8'h72,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* XOR,C,A */
                {8'h82,8'hxx,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* INC,,C */
                {8'h92,8'hxx,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* DEC,,C */
                {8'ha3,8'hxx,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* INCW,,BC */
                {8'hb3,8'hxx,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* DECW,,BC */
                {8'h31,8'h07,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHL,C,0 */
                {8'h31,8'h17,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHL,C,1 */
                {8'h31,8'h27,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHL,C,2 */
                {8'h31,8'h37,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHL,C,3 */
                {8'h31,8'h47,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHL,C,4 */
                {8'h31,8'h57,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHL,C,5 */
                {8'h31,8'h67,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHL,C,6 */
                {8'h31,8'h77,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHL,C,7 */
                {8'h31,8'h0c,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHLW,BC,0 */
                {8'h31,8'h1c,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHLW,BC,1 */
                {8'h31,8'h2c,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHLW,BC,2 */
                {8'h31,8'h3c,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHLW,BC,3 */
                {8'h31,8'h4c,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHLW,BC,4 */
                {8'h31,8'h5c,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHLW,BC,5 */
                {8'h31,8'h6c,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHLW,BC,6 */
                {8'h31,8'h7c,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHLW,BC,7 */
                {8'h31,8'h8c,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHLW,BC,8 */
                {8'h31,8'h9c,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHLW,BC,9 */
                {8'h31,8'hac,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHLW,BC,10 */
                {8'h31,8'hbc,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHLW,BC,11 */
                {8'h31,8'hcc,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHLW,BC,12 */
                {8'h31,8'hdc,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHLW,BC,13 */
                {8'h31,8'hec,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHLW,BC,14 */
                {8'h31,8'hfc,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHLW,BC,15 */
                {8'h61,8'hfe,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* ROLWC,BC,1 */
                {8'hc2,8'hxx,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* POP,,BC */
                {8'h61,8'h9a,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* XCH,A,C */
                {8'h31,8'h87,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHL,C,0 */
                {8'h31,8'h97,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHL,C,1 */
                {8'h31,8'ha7,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHL,C,2 */
                {8'h31,8'hb7,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHL,C,3 */
                {8'h31,8'hc7,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHL,C,4 */
                {8'h31,8'hd7,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHL,C,5 */
                {8'h31,8'he7,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHL,C,6 */
                {8'h31,8'hf7,2'bxx} : dec_C_enable_adrstage = 1'b1;  /* SHL,C,7 */
                default : dec_C_enable_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_C_enable <= 1'b0;
        else if(cpuen) dec_C_enable <= dec_C_enable_adrstage;
    end
    output dec_D_enable;
    reg    dec_D_enable, dec_D_enable_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1|| skpack == 1'b1) begin
            dec_D_enable_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h55,8'hxx,2'bxx} : dec_D_enable_adrstage = 1'b1;  /* MOV,D,#byte */
                {8'h75,8'hxx,2'bxx} : dec_D_enable_adrstage = 1'b1;  /* MOV,D,A */
                {8'h61,8'h8d,2'bxx} : dec_D_enable_adrstage = 1'b1;  /* XCH,A,D */
                {8'h34,8'hxx,2'bxx} : dec_D_enable_adrstage = 1'b1;  /* MOVW,DE,#word */
                {8'h14,8'hxx,2'bxx} : dec_D_enable_adrstage = 1'b1;  /* MOVW,DE,AX */
                {8'hea,8'hxx,2'bxx} : dec_D_enable_adrstage = 1'b1;  /* MOVW,DE,saddrp */
                {8'heb,8'hxx,2'bxx} : dec_D_enable_adrstage = 1'b1;  /* MOVW,DE,!addr16 */
                {8'h35,8'hxx,2'bxx} : dec_D_enable_adrstage = 1'b1;  /* XCHW,AX,DE */
                {8'h61,8'h05,2'bxx} : dec_D_enable_adrstage = 1'b1;  /* ADD,D,A */
                {8'h61,8'h15,2'bxx} : dec_D_enable_adrstage = 1'b1;  /* ADDC,D,A */
                {8'h61,8'h25,2'bxx} : dec_D_enable_adrstage = 1'b1;  /* SUB,D,A */
                {8'h61,8'h35,2'bxx} : dec_D_enable_adrstage = 1'b1;  /* SUBC,D,A */
                {8'h61,8'h55,2'bxx} : dec_D_enable_adrstage = 1'b1;  /* AND,D,A */
                {8'h61,8'h65,2'bxx} : dec_D_enable_adrstage = 1'b1;  /* OR,D,A */
                {8'h61,8'h75,2'bxx} : dec_D_enable_adrstage = 1'b1;  /* XOR,D,A */
                {8'h85,8'hxx,2'bxx} : dec_D_enable_adrstage = 1'b1;  /* INC,,D */
                {8'h95,8'hxx,2'bxx} : dec_D_enable_adrstage = 1'b1;  /* DEC,,D */
                {8'ha5,8'hxx,2'bxx} : dec_D_enable_adrstage = 1'b1;  /* INCW,,DE */
                {8'hb5,8'hxx,2'bxx} : dec_D_enable_adrstage = 1'b1;  /* DECW,,DE */
                {8'hc4,8'hxx,2'bxx} : dec_D_enable_adrstage = 1'b1;  /* POP,,DE */
                {8'h61,8'h9d,2'bxx} : dec_D_enable_adrstage = 1'b1;  /* XCH,A,D */
                default : dec_D_enable_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_D_enable <= 1'b0;
        else if(cpuen) dec_D_enable <= dec_D_enable_adrstage;
    end
    output dec_E_enable;
    reg    dec_E_enable, dec_E_enable_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1|| skpack == 1'b1) begin
            dec_E_enable_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h54,8'hxx,2'bxx} : dec_E_enable_adrstage = 1'b1;  /* MOV,E,#byte */
                {8'h74,8'hxx,2'bxx} : dec_E_enable_adrstage = 1'b1;  /* MOV,E,A */
                {8'h61,8'h8c,2'bxx} : dec_E_enable_adrstage = 1'b1;  /* XCH,A,E */
                {8'h34,8'hxx,2'bxx} : dec_E_enable_adrstage = 1'b1;  /* MOVW,DE,#word */
                {8'h14,8'hxx,2'bxx} : dec_E_enable_adrstage = 1'b1;  /* MOVW,DE,AX */
                {8'hea,8'hxx,2'bxx} : dec_E_enable_adrstage = 1'b1;  /* MOVW,DE,saddrp */
                {8'heb,8'hxx,2'bxx} : dec_E_enable_adrstage = 1'b1;  /* MOVW,DE,!addr16 */
                {8'h35,8'hxx,2'bxx} : dec_E_enable_adrstage = 1'b1;  /* XCHW,AX,DE */
                {8'h61,8'h04,2'bxx} : dec_E_enable_adrstage = 1'b1;  /* ADD,E,A */
                {8'h61,8'h14,2'bxx} : dec_E_enable_adrstage = 1'b1;  /* ADDC,E,A */
                {8'h61,8'h24,2'bxx} : dec_E_enable_adrstage = 1'b1;  /* SUB,E,A */
                {8'h61,8'h34,2'bxx} : dec_E_enable_adrstage = 1'b1;  /* SUBC,E,A */
                {8'h61,8'h54,2'bxx} : dec_E_enable_adrstage = 1'b1;  /* AND,E,A */
                {8'h61,8'h64,2'bxx} : dec_E_enable_adrstage = 1'b1;  /* OR,E,A */
                {8'h61,8'h74,2'bxx} : dec_E_enable_adrstage = 1'b1;  /* XOR,E,A */
                {8'h84,8'hxx,2'bxx} : dec_E_enable_adrstage = 1'b1;  /* INC,,E */
                {8'h94,8'hxx,2'bxx} : dec_E_enable_adrstage = 1'b1;  /* DEC,,E */
                {8'ha5,8'hxx,2'bxx} : dec_E_enable_adrstage = 1'b1;  /* INCW,,DE */
                {8'hb5,8'hxx,2'bxx} : dec_E_enable_adrstage = 1'b1;  /* DECW,,DE */
                {8'hc4,8'hxx,2'bxx} : dec_E_enable_adrstage = 1'b1;  /* POP,,DE */
                {8'h61,8'h9c,2'bxx} : dec_E_enable_adrstage = 1'b1;  /* XCH,A,E */
                default : dec_E_enable_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_E_enable <= 1'b0;
        else if(cpuen) dec_E_enable <= dec_E_enable_adrstage;
    end
    output dec_H_enable;
    reg    dec_H_enable, dec_H_enable_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1|| skpack == 1'b1) begin
            dec_H_enable_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h57,8'hxx,2'bxx} : dec_H_enable_adrstage = 1'b1;  /* MOV,H,#byte */
                {8'h77,8'hxx,2'bxx} : dec_H_enable_adrstage = 1'b1;  /* MOV,H,A */
                {8'h61,8'h8f,2'bxx} : dec_H_enable_adrstage = 1'b1;  /* XCH,A,H */
                {8'h36,8'hxx,2'bxx} : dec_H_enable_adrstage = 1'b1;  /* MOVW,HL,#word */
                {8'h16,8'hxx,2'bxx} : dec_H_enable_adrstage = 1'b1;  /* MOVW,HL,AX */
                {8'hfa,8'hxx,2'bxx} : dec_H_enable_adrstage = 1'b1;  /* MOVW,HL,saddrp */
                {8'hfb,8'hxx,2'bxx} : dec_H_enable_adrstage = 1'b1;  /* MOVW,HL,!addr16 */
                {8'h37,8'hxx,2'bxx} : dec_H_enable_adrstage = 1'b1;  /* XCHW,AX,HL */
                {8'h61,8'h07,2'bxx} : dec_H_enable_adrstage = 1'b1;  /* ADD,H,A */
                {8'h61,8'h17,2'bxx} : dec_H_enable_adrstage = 1'b1;  /* ADDC,H,A */
                {8'h61,8'h27,2'bxx} : dec_H_enable_adrstage = 1'b1;  /* SUB,H,A */
                {8'h61,8'h37,2'bxx} : dec_H_enable_adrstage = 1'b1;  /* SUBC,H,A */
                {8'h61,8'h57,2'bxx} : dec_H_enable_adrstage = 1'b1;  /* AND,H,A */
                {8'h61,8'h67,2'bxx} : dec_H_enable_adrstage = 1'b1;  /* OR,H,A */
                {8'h61,8'h77,2'bxx} : dec_H_enable_adrstage = 1'b1;  /* XOR,H,A */
                {8'h87,8'hxx,2'bxx} : dec_H_enable_adrstage = 1'b1;  /* INC,,H */
                {8'h97,8'hxx,2'bxx} : dec_H_enable_adrstage = 1'b1;  /* DEC,,H */
                {8'ha7,8'hxx,2'bxx} : dec_H_enable_adrstage = 1'b1;  /* INCW,,HL */
                {8'hb7,8'hxx,2'bxx} : dec_H_enable_adrstage = 1'b1;  /* DECW,,HL */
                {8'hc6,8'hxx,2'bxx} : dec_H_enable_adrstage = 1'b1;  /* POP,,HL */
                {8'h61,8'h9f,2'bxx} : dec_H_enable_adrstage = 1'b1;  /* XCH,A,H */
                default : dec_H_enable_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_H_enable <= 1'b0;
        else if(cpuen) dec_H_enable <= dec_H_enable_adrstage;
    end
    output dec_L_enable;
    reg    dec_L_enable, dec_L_enable_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1|| skpack == 1'b1) begin
            dec_L_enable_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h56,8'hxx,2'bxx} : dec_L_enable_adrstage = 1'b1;  /* MOV,L,#byte */
                {8'h76,8'hxx,2'bxx} : dec_L_enable_adrstage = 1'b1;  /* MOV,L,A */
                {8'h61,8'h8e,2'bxx} : dec_L_enable_adrstage = 1'b1;  /* XCH,A,L */
                {8'h36,8'hxx,2'bxx} : dec_L_enable_adrstage = 1'b1;  /* MOVW,HL,#word */
                {8'h16,8'hxx,2'bxx} : dec_L_enable_adrstage = 1'b1;  /* MOVW,HL,AX */
                {8'hfa,8'hxx,2'bxx} : dec_L_enable_adrstage = 1'b1;  /* MOVW,HL,saddrp */
                {8'hfb,8'hxx,2'bxx} : dec_L_enable_adrstage = 1'b1;  /* MOVW,HL,!addr16 */
                {8'h37,8'hxx,2'bxx} : dec_L_enable_adrstage = 1'b1;  /* XCHW,AX,HL */
                {8'h61,8'h06,2'bxx} : dec_L_enable_adrstage = 1'b1;  /* ADD,L,A */
                {8'h61,8'h16,2'bxx} : dec_L_enable_adrstage = 1'b1;  /* ADDC,L,A */
                {8'h61,8'h26,2'bxx} : dec_L_enable_adrstage = 1'b1;  /* SUB,L,A */
                {8'h61,8'h36,2'bxx} : dec_L_enable_adrstage = 1'b1;  /* SUBC,L,A */
                {8'h61,8'h56,2'bxx} : dec_L_enable_adrstage = 1'b1;  /* AND,L,A */
                {8'h61,8'h66,2'bxx} : dec_L_enable_adrstage = 1'b1;  /* OR,L,A */
                {8'h61,8'h76,2'bxx} : dec_L_enable_adrstage = 1'b1;  /* XOR,L,A */
                {8'h86,8'hxx,2'bxx} : dec_L_enable_adrstage = 1'b1;  /* INC,,L */
                {8'h96,8'hxx,2'bxx} : dec_L_enable_adrstage = 1'b1;  /* DEC,,L */
                {8'ha7,8'hxx,2'bxx} : dec_L_enable_adrstage = 1'b1;  /* INCW,,HL */
                {8'hb7,8'hxx,2'bxx} : dec_L_enable_adrstage = 1'b1;  /* DECW,,HL */
                {8'hc6,8'hxx,2'bxx} : dec_L_enable_adrstage = 1'b1;  /* POP,,HL */
                {8'h61,8'h9e,2'bxx} : dec_L_enable_adrstage = 1'b1;  /* XCH,A,L */
                default : dec_L_enable_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_L_enable <= 1'b0;
        else if(cpuen) dec_L_enable <= dec_L_enable_adrstage;
    end
    output dec_ES_enable;
    reg    dec_ES_enable, dec_ES_enable_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1|| skpack == 1'b1) begin
            dec_ES_enable_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h41,8'hxx,2'bxx} : dec_ES_enable_adrstage = 1'b1;  /* MOV,ES,#byte */
                {8'h61,8'hb8,2'bxx} : dec_ES_enable_adrstage = 1'b1;  /* MOV,ES,saddr */
                default : dec_ES_enable_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_ES_enable <= 1'b0;
        else if(cpuen) dec_ES_enable <= dec_ES_enable_adrstage;
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*����ADD,ADDC,SUB,SUBC,AND,OR,XOR,INC,DEC��					*/
/*���������������ꥢ�������黻�򣲥���å��ܤ��飱����å��ܤ��ѹ�		*/
/*------------------------------------------------------------------------------*/

    output dec_Z_enable;
    reg    dec_Z_enable, dec_Z_enable_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1|| skpack == 1'b1) begin
            dec_Z_enable_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h0c,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,A,#byte */
                {8'h0a,8'hxx,2'bx0} : dec_Z_enable_adrstage = 1'b1;  /* ADD,saddr,#byte */
                {8'h61,8'h08,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,A,X */
                {8'h61,8'h0a,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,A,C */
                {8'h61,8'h0b,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,A,B */
                {8'h61,8'h0c,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,A,E */
                {8'h61,8'h0d,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,A,D */
                {8'h61,8'h0e,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,A,L */
                {8'h61,8'h0f,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,A,H */
                {8'h61,8'h00,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,X,A */
                {8'h61,8'h01,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,A,A */
                {8'h61,8'h02,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,C,A */
                {8'h61,8'h03,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,B,A */
                {8'h61,8'h04,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,E,A */
                {8'h61,8'h05,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,D,A */
                {8'h61,8'h06,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,L,A */
                {8'h61,8'h07,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,H,A */
                {8'h0b,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,A,saddr */
                {8'h0f,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,A,!addr16 */
                {8'h0d,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,A,[HL] */
                {8'h0e,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,A,[HL+byte] */
                {8'h61,8'h80,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,A,[HL+B] */
                {8'h61,8'h82,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,A,[HL+C] */
                {8'h1c,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,A,#byte */
                {8'h1a,8'hxx,2'bx0} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,saddr,#byte */
                {8'h61,8'h18,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,A,X */
                {8'h61,8'h1a,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,A,C */
                {8'h61,8'h1b,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,A,B */
                {8'h61,8'h1c,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,A,E */
                {8'h61,8'h1d,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,A,D */
                {8'h61,8'h1e,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,A,L */
                {8'h61,8'h1f,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,A,H */
                {8'h61,8'h10,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,X,A */
                {8'h61,8'h11,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,A,A */
                {8'h61,8'h12,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,C,A */
                {8'h61,8'h13,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,B,A */
                {8'h61,8'h14,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,E,A */
                {8'h61,8'h15,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,D,A */
                {8'h61,8'h16,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,L,A */
                {8'h61,8'h17,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,H,A */
                {8'h1b,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,A,saddr */
                {8'h1f,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,A,!addr16 */
                {8'h1d,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,A,[HL] */
                {8'h1e,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,A,[HL+byte] */
                {8'h61,8'h90,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,A,[HL+B] */
                {8'h61,8'h92,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,A,[HL+C] */
                {8'h2c,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,A,#byte */
                {8'h2a,8'hxx,2'bx0} : dec_Z_enable_adrstage = 1'b1;  /* SUB,saddr,#byte */
                {8'h61,8'h28,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,A,X */
                {8'h61,8'h2a,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,A,C */
                {8'h61,8'h2b,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,A,B */
                {8'h61,8'h2c,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,A,E */
                {8'h61,8'h2d,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,A,D */
                {8'h61,8'h2e,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,A,L */
                {8'h61,8'h2f,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,A,H */
                {8'h61,8'h20,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,X,A */
                {8'h61,8'h21,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,A,A */
                {8'h61,8'h22,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,C,A */
                {8'h61,8'h23,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,B,A */
                {8'h61,8'h24,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,E,A */
                {8'h61,8'h25,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,D,A */
                {8'h61,8'h26,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,L,A */
                {8'h61,8'h27,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,H,A */
                {8'h2b,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,A,saddr */
                {8'h2f,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,A,!addr16 */
                {8'h2d,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,A,[HL] */
                {8'h2e,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,A,[HL+byte] */
                {8'h61,8'ha0,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,A,[HL+B] */
                {8'h61,8'ha2,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,A,[HL+C] */
                {8'h3c,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,A,#byte */
                {8'h3a,8'hxx,2'bx0} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,saddr,#byte */
                {8'h61,8'h38,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,A,X */
                {8'h61,8'h3a,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,A,C */
                {8'h61,8'h3b,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,A,B */
                {8'h61,8'h3c,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,A,E */
                {8'h61,8'h3d,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,A,D */
                {8'h61,8'h3e,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,A,L */
                {8'h61,8'h3f,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,A,H */
                {8'h61,8'h30,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,X,A */
                {8'h61,8'h31,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,A,A */
                {8'h61,8'h32,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,C,A */
                {8'h61,8'h33,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,B,A */
                {8'h61,8'h34,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,E,A */
                {8'h61,8'h35,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,D,A */
                {8'h61,8'h36,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,L,A */
                {8'h61,8'h37,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,H,A */
                {8'h3b,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,A,saddr */
                {8'h3f,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,A,!addr16 */
                {8'h3d,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,A,[HL] */
                {8'h3e,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,A,[HL+byte] */
                {8'h61,8'hb0,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,A,[HL+B] */
                {8'h61,8'hb2,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,A,[HL+C] */
                {8'h5c,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,A,#byte */
                {8'h5a,8'hxx,2'bx0} : dec_Z_enable_adrstage = 1'b1;  /* AND,saddr,#byte */
                {8'h61,8'h58,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,A,X */
                {8'h61,8'h5a,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,A,C */
                {8'h61,8'h5b,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,A,B */
                {8'h61,8'h5c,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,A,E */
                {8'h61,8'h5d,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,A,D */
                {8'h61,8'h5e,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,A,L */
                {8'h61,8'h5f,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,A,H */
                {8'h61,8'h50,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,X,A */
                {8'h61,8'h51,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,A,A */
                {8'h61,8'h52,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,C,A */
                {8'h61,8'h53,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,B,A */
                {8'h61,8'h54,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,E,A */
                {8'h61,8'h55,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,D,A */
                {8'h61,8'h56,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,L,A */
                {8'h61,8'h57,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,H,A */
                {8'h5b,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,A,saddr */
                {8'h5f,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,A,!addr16 */
                {8'h5d,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,A,[HL] */
                {8'h5e,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,A,[HL+byte] */
                {8'h61,8'hd0,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,A,[HL+B] */
                {8'h61,8'hd2,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,A,[HL+C] */
                {8'h6c,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,A,#byte */
                {8'h6a,8'hxx,2'bx0} : dec_Z_enable_adrstage = 1'b1;  /* OR,saddr,#byte */
                {8'h61,8'h68,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,A,X */
                {8'h61,8'h6a,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,A,C */
                {8'h61,8'h6b,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,A,B */
                {8'h61,8'h6c,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,A,E */
                {8'h61,8'h6d,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,A,D */
                {8'h61,8'h6e,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,A,L */
                {8'h61,8'h6f,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,A,H */
                {8'h61,8'h60,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,X,A */
                {8'h61,8'h61,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,A,A */
                {8'h61,8'h62,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,C,A */
                {8'h61,8'h63,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,B,A */
                {8'h61,8'h64,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,E,A */
                {8'h61,8'h65,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,D,A */
                {8'h61,8'h66,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,L,A */
                {8'h61,8'h67,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,H,A */
                {8'h6b,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,A,saddr */
                {8'h6f,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,A,!addr16 */
                {8'h6d,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,A,[HL] */
                {8'h6e,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,A,[HL+byte] */
                {8'h61,8'he0,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,A,[HL+B] */
                {8'h61,8'he2,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,A,[HL+C] */
                {8'h7c,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,A,#byte */
                {8'h7a,8'hxx,2'bx0} : dec_Z_enable_adrstage = 1'b1;  /* XOR,saddr,#byte */
                {8'h61,8'h78,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,A,X */
                {8'h61,8'h7a,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,A,C */
                {8'h61,8'h7b,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,A,B */
                {8'h61,8'h7c,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,A,E */
                {8'h61,8'h7d,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,A,D */
                {8'h61,8'h7e,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,A,L */
                {8'h61,8'h7f,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,A,H */
                {8'h61,8'h70,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,X,A */
                {8'h61,8'h71,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,A,A */
                {8'h61,8'h72,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,C,A */
                {8'h61,8'h73,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,B,A */
                {8'h61,8'h74,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,E,A */
                {8'h61,8'h75,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,D,A */
                {8'h61,8'h76,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,L,A */
                {8'h61,8'h77,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,H,A */
                {8'h7b,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,A,saddr */
                {8'h7f,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,A,!addr16 */
                {8'h7d,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,A,[HL] */
                {8'h7e,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,A,[HL+byte] */
                {8'h61,8'hf0,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,A,[HL+B] */
                {8'h61,8'hf2,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,A,[HL+C] */
                {8'h4c,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,A,#byte */
                {8'h4a,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,saddr,#byte */
                {8'h40,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,!addr16,#byte */
                {8'h61,8'h48,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,A,X */
                {8'h61,8'h4a,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,A,C */
                {8'h61,8'h4b,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,A,B */
                {8'h61,8'h4c,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,A,E */
                {8'h61,8'h4d,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,A,D */
                {8'h61,8'h4e,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,A,L */
                {8'h61,8'h4f,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,A,H */
                {8'h61,8'h40,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,X,A */
                {8'h61,8'h41,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,A,A */
                {8'h61,8'h42,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,C,A */
                {8'h61,8'h43,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,B,A */
                {8'h61,8'h44,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,E,A */
                {8'h61,8'h45,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,D,A */
                {8'h61,8'h46,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,L,A */
                {8'h61,8'h47,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,H,A */
                {8'h4b,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,A,saddr */
                {8'h4f,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,A,!addr16 */
                {8'h4d,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,A,[HL] */
                {8'h4e,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,A,[HL+byte] */
                {8'h61,8'hc0,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,A,[HL+B] */
                {8'h61,8'hc2,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP,A,[HL+C] */
                {8'h61,8'hde,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMPS,X,[HL+byte] */
                {8'hd1,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP0,,A */
                {8'hd0,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP0,,X */
                {8'hd3,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP0,,B */
                {8'hd2,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP0,,C */
                {8'hd4,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP0,,saddr */
                {8'hd5,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMP0,,!addr16 */
                {8'h04,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDW,AX,#word */
                {8'h01,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDW,AX,AX */
                {8'h03,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDW,AX,BC */
                {8'h05,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDW,AX,DE */
                {8'h07,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDW,AX,HL */
                {8'h06,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDW,AX,saddrp */
                {8'h02,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDW,AX,!addr16 */
                {8'h61,8'h09,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDW,AX,[HL+byte] */
                {8'h24,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBW,AX,#word */
                {8'h21,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBW,AX,AX */
                {8'h23,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBW,AX,BC */
                {8'h25,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBW,AX,DE */
                {8'h27,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBW,AX,HL */
                {8'h26,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBW,AX,saddrp */
                {8'h22,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBW,AX,!addr16 */
                {8'h61,8'h29,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBW,AX,[HL+byte] */
                {8'h44,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMPW,AX,#word */
                {8'h43,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMPW,AX,BC */
                {8'h45,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMPW,AX,DE */
                {8'h47,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMPW,AX,HL */
                {8'h46,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMPW,AX,saddrp */
                {8'h42,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMPW,AX,!addr16 */
                {8'h61,8'h49,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* CMPW,AX,[HL+byte] */
                {8'h80,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* INC,,X */
                {8'h81,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* INC,,A */
                {8'h82,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* INC,,C */
                {8'h83,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* INC,,B */
                {8'h84,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* INC,,E */
                {8'h85,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* INC,,D */
                {8'h86,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* INC,,L */
                {8'h87,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* INC,,H */
                {8'ha4,8'hxx,2'bx0} : dec_Z_enable_adrstage = 1'b1;  /* INC,,saddr */
                {8'ha0,8'hxx,2'bx0} : dec_Z_enable_adrstage = 1'b1;  /* INC,,!addr16 */
                {8'h61,8'h59,2'bx0} : dec_Z_enable_adrstage = 1'b1;  /* INC,,[HL+byte] */
                {8'h90,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* DEC,,X */
                {8'h91,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* DEC,,A */
                {8'h92,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* DEC,,C */
                {8'h93,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* DEC,,B */
                {8'h94,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* DEC,,E */
                {8'h95,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* DEC,,D */
                {8'h96,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* DEC,,L */
                {8'h97,8'hxx,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* DEC,,H */
                {8'hb4,8'hxx,2'bx0} : dec_Z_enable_adrstage = 1'b1;  /* DEC,,saddr */
                {8'hb0,8'hxx,2'bx0} : dec_Z_enable_adrstage = 1'b1;  /* DEC,,!addr16 */
                {8'h61,8'h69,2'bx0} : dec_Z_enable_adrstage = 1'b1;  /* DEC,,[HL+byte] */
                {8'h61,8'hec,2'b01} : dec_Z_enable_adrstage = 1'b1;  /* RETB,, */
                {8'h61,8'hfc,2'b01} : dec_Z_enable_adrstage = 1'b1;  /* RETI,, */
                {8'h61,8'hcd,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* POP,,PSW */
                {8'h61,8'h19,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,A,A */
                {8'h61,8'h39,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,A,A */
                {8'h61,8'hd1,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* AND,A,[HL+B] */
                {8'h61,8'he1,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* OR,A,[HL+B] */
                {8'h61,8'hf1,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* XOR,A,[HL+B] */
                {8'h61,8'h83,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADD,A,[HL+C] */
                {8'h61,8'h93,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* ADDC,A,[HL+C] */
                {8'h61,8'ha3,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUB,A,[HL+C] */
                {8'h61,8'hb3,2'bxx} : dec_Z_enable_adrstage = 1'b1;  /* SUBC,A,[HL+C] */
                default : dec_Z_enable_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_Z_enable <= 1'b0;
        else if(cpuen) dec_Z_enable <= dec_Z_enable_adrstage;
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*����ADD,ADDC,SUB,SUBC��							*/
/*���������������ꥢ�������黻�򣲥���å��ܤ��飱����å��ܤ��ѹ�		*/
/*------------------------------------------------------------------------------*/

    output dec_CY_enable;
    reg    dec_CY_enable, dec_CY_enable_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1|| skpack == 1'b1) begin
            dec_CY_enable_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h0c,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,A,#byte */
                {8'h0a,8'hxx,2'bx0} : dec_CY_enable_adrstage = 1'b1;  /* ADD,saddr,#byte */
                {8'h61,8'h08,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,A,X */
                {8'h61,8'h0a,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,A,C */
                {8'h61,8'h0b,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,A,B */
                {8'h61,8'h0c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,A,E */
                {8'h61,8'h0d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,A,D */
                {8'h61,8'h0e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,A,L */
                {8'h61,8'h0f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,A,H */
                {8'h61,8'h00,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,X,A */
                {8'h61,8'h01,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,A,A */
                {8'h61,8'h02,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,C,A */
                {8'h61,8'h03,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,B,A */
                {8'h61,8'h04,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,E,A */
                {8'h61,8'h05,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,D,A */
                {8'h61,8'h06,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,L,A */
                {8'h61,8'h07,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,H,A */
                {8'h0b,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,A,saddr */
                {8'h0f,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,A,!addr16 */
                {8'h0d,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,A,[HL] */
                {8'h0e,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,A,[HL+byte] */
                {8'h61,8'h80,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,A,[HL+B] */
                {8'h61,8'h82,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,A,[HL+C] */
                {8'h1c,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,A,#byte */
                {8'h1a,8'hxx,2'bx0} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,saddr,#byte */
                {8'h61,8'h18,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,A,X */
                {8'h61,8'h1a,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,A,C */
                {8'h61,8'h1b,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,A,B */
                {8'h61,8'h1c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,A,E */
                {8'h61,8'h1d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,A,D */
                {8'h61,8'h1e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,A,L */
                {8'h61,8'h1f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,A,H */
                {8'h61,8'h10,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,X,A */
                {8'h61,8'h11,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,A,A */
                {8'h61,8'h12,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,C,A */
                {8'h61,8'h13,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,B,A */
                {8'h61,8'h14,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,E,A */
                {8'h61,8'h15,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,D,A */
                {8'h61,8'h16,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,L,A */
                {8'h61,8'h17,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,H,A */
                {8'h1b,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,A,saddr */
                {8'h1f,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,A,!addr16 */
                {8'h1d,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,A,[HL] */
                {8'h1e,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,A,[HL+byte] */
                {8'h61,8'h90,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,A,[HL+B] */
                {8'h61,8'h92,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,A,[HL+C] */
                {8'h2c,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,A,#byte */
                {8'h2a,8'hxx,2'bx0} : dec_CY_enable_adrstage = 1'b1;  /* SUB,saddr,#byte */
                {8'h61,8'h28,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,A,X */
                {8'h61,8'h2a,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,A,C */
                {8'h61,8'h2b,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,A,B */
                {8'h61,8'h2c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,A,E */
                {8'h61,8'h2d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,A,D */
                {8'h61,8'h2e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,A,L */
                {8'h61,8'h2f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,A,H */
                {8'h61,8'h20,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,X,A */
                {8'h61,8'h21,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,A,A */
                {8'h61,8'h22,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,C,A */
                {8'h61,8'h23,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,B,A */
                {8'h61,8'h24,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,E,A */
                {8'h61,8'h25,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,D,A */
                {8'h61,8'h26,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,L,A */
                {8'h61,8'h27,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,H,A */
                {8'h2b,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,A,saddr */
                {8'h2f,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,A,!addr16 */
                {8'h2d,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,A,[HL] */
                {8'h2e,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,A,[HL+byte] */
                {8'h61,8'ha0,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,A,[HL+B] */
                {8'h61,8'ha2,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,A,[HL+C] */
                {8'h3c,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,A,#byte */
                {8'h3a,8'hxx,2'bx0} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,saddr,#byte */
                {8'h61,8'h38,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,A,X */
                {8'h61,8'h3a,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,A,C */
                {8'h61,8'h3b,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,A,B */
                {8'h61,8'h3c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,A,E */
                {8'h61,8'h3d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,A,D */
                {8'h61,8'h3e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,A,L */
                {8'h61,8'h3f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,A,H */
                {8'h61,8'h30,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,X,A */
                {8'h61,8'h31,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,A,A */
                {8'h61,8'h32,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,C,A */
                {8'h61,8'h33,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,B,A */
                {8'h61,8'h34,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,E,A */
                {8'h61,8'h35,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,D,A */
                {8'h61,8'h36,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,L,A */
                {8'h61,8'h37,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,H,A */
                {8'h3b,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,A,saddr */
                {8'h3f,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,A,!addr16 */
                {8'h3d,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,A,[HL] */
                {8'h3e,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,A,[HL+byte] */
                {8'h61,8'hb0,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,A,[HL+B] */
                {8'h61,8'hb2,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,A,[HL+C] */
                {8'h4c,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,A,#byte */
                {8'h4a,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,saddr,#byte */
                {8'h40,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,!addr16,#byte */
                {8'h61,8'h48,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,A,X */
                {8'h61,8'h4a,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,A,C */
                {8'h61,8'h4b,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,A,B */
                {8'h61,8'h4c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,A,E */
                {8'h61,8'h4d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,A,D */
                {8'h61,8'h4e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,A,L */
                {8'h61,8'h4f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,A,H */
                {8'h61,8'h40,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,X,A */
                {8'h61,8'h41,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,A,A */
                {8'h61,8'h42,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,C,A */
                {8'h61,8'h43,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,B,A */
                {8'h61,8'h44,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,E,A */
                {8'h61,8'h45,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,D,A */
                {8'h61,8'h46,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,L,A */
                {8'h61,8'h47,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,H,A */
                {8'h4b,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,A,saddr */
                {8'h4f,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,A,!addr16 */
                {8'h4d,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,A,[HL] */
                {8'h4e,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,A,[HL+byte] */
                {8'h61,8'hc0,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,A,[HL+B] */
                {8'h61,8'hc2,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP,A,[HL+C] */
                {8'h61,8'hde,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMPS,X,[HL+byte] */
                {8'hd1,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP0,,A */
                {8'hd0,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP0,,X */
                {8'hd3,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP0,,B */
                {8'hd2,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP0,,C */
                {8'hd4,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP0,,saddr */
                {8'hd5,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMP0,,!addr16 */
                {8'h04,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDW,AX,#word */
                {8'h01,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDW,AX,AX */
                {8'h03,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDW,AX,BC */
                {8'h05,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDW,AX,DE */
                {8'h07,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDW,AX,HL */
                {8'h06,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDW,AX,saddrp */
                {8'h02,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDW,AX,!addr16 */
                {8'h61,8'h09,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDW,AX,[HL+byte] */
                {8'h24,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBW,AX,#word */
                {8'h21,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBW,AX,AX */
                {8'h23,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBW,AX,BC */
                {8'h25,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBW,AX,DE */
                {8'h27,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBW,AX,HL */
                {8'h26,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBW,AX,saddrp */
                {8'h22,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBW,AX,!addr16 */
                {8'h61,8'h29,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBW,AX,[HL+byte] */
                {8'h44,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMPW,AX,#word */
                {8'h43,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMPW,AX,BC */
                {8'h45,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMPW,AX,DE */
                {8'h47,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMPW,AX,HL */
                {8'h46,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMPW,AX,saddrp */
                {8'h42,8'hxx,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMPW,AX,!addr16 */
                {8'h61,8'h49,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CMPW,AX,[HL+byte] */
                {8'h31,8'h0a,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHR,A,0 */
                {8'h31,8'h1a,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHR,A,1 */
                {8'h31,8'h2a,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHR,A,2 */
                {8'h31,8'h3a,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHR,A,3 */
                {8'h31,8'h4a,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHR,A,4 */
                {8'h31,8'h5a,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHR,A,5 */
                {8'h31,8'h6a,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHR,A,6 */
                {8'h31,8'h7a,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHR,A,7 */
                {8'h31,8'h0e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHRW,AX,0 */
                {8'h31,8'h1e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHRW,AX,1 */
                {8'h31,8'h2e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHRW,AX,2 */
                {8'h31,8'h3e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHRW,AX,3 */
                {8'h31,8'h4e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHRW,AX,4 */
                {8'h31,8'h5e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHRW,AX,5 */
                {8'h31,8'h6e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHRW,AX,6 */
                {8'h31,8'h7e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHRW,AX,7 */
                {8'h31,8'h8e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHRW,AX,8 */
                {8'h31,8'h9e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHRW,AX,9 */
                {8'h31,8'hae,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHRW,AX,10 */
                {8'h31,8'hbe,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHRW,AX,11 */
                {8'h31,8'hce,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHRW,AX,12 */
                {8'h31,8'hde,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHRW,AX,13 */
                {8'h31,8'hee,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHRW,AX,14 */
                {8'h31,8'hfe,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHRW,AX,15 */
                {8'h31,8'h09,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,A,0 */
                {8'h31,8'h19,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,A,1 */
                {8'h31,8'h29,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,A,2 */
                {8'h31,8'h39,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,A,3 */
                {8'h31,8'h49,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,A,4 */
                {8'h31,8'h59,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,A,5 */
                {8'h31,8'h69,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,A,6 */
                {8'h31,8'h79,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,A,7 */
                {8'h31,8'h08,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,B,0 */
                {8'h31,8'h18,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,B,1 */
                {8'h31,8'h28,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,B,2 */
                {8'h31,8'h38,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,B,3 */
                {8'h31,8'h48,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,B,4 */
                {8'h31,8'h58,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,B,5 */
                {8'h31,8'h68,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,B,6 */
                {8'h31,8'h78,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,B,7 */
                {8'h31,8'h07,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,C,0 */
                {8'h31,8'h17,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,C,1 */
                {8'h31,8'h27,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,C,2 */
                {8'h31,8'h37,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,C,3 */
                {8'h31,8'h47,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,C,4 */
                {8'h31,8'h57,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,C,5 */
                {8'h31,8'h67,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,C,6 */
                {8'h31,8'h77,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,C,7 */
                {8'h31,8'h0d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,AX,0 */
                {8'h31,8'h1d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,AX,1 */
                {8'h31,8'h2d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,AX,2 */
                {8'h31,8'h3d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,AX,3 */
                {8'h31,8'h4d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,AX,4 */
                {8'h31,8'h5d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,AX,5 */
                {8'h31,8'h6d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,AX,6 */
                {8'h31,8'h7d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,AX,7 */
                {8'h31,8'h8d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,AX,8 */
                {8'h31,8'h9d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,AX,9 */
                {8'h31,8'had,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,AX,10 */
                {8'h31,8'hbd,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,AX,11 */
                {8'h31,8'hcd,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,AX,12 */
                {8'h31,8'hdd,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,AX,13 */
                {8'h31,8'hed,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,AX,14 */
                {8'h31,8'hfd,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,AX,15 */
                {8'h31,8'h0c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,BC,0 */
                {8'h31,8'h1c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,BC,1 */
                {8'h31,8'h2c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,BC,2 */
                {8'h31,8'h3c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,BC,3 */
                {8'h31,8'h4c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,BC,4 */
                {8'h31,8'h5c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,BC,5 */
                {8'h31,8'h6c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,BC,6 */
                {8'h31,8'h7c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,BC,7 */
                {8'h31,8'h8c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,BC,8 */
                {8'h31,8'h9c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,BC,9 */
                {8'h31,8'hac,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,BC,10 */
                {8'h31,8'hbc,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,BC,11 */
                {8'h31,8'hcc,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,BC,12 */
                {8'h31,8'hdc,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,BC,13 */
                {8'h31,8'hec,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,BC,14 */
                {8'h31,8'hfc,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHLW,BC,15 */
                {8'h31,8'h0b,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SAR,A,0 */
                {8'h31,8'h1b,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SAR,A,1 */
                {8'h31,8'h2b,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SAR,A,2 */
                {8'h31,8'h3b,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SAR,A,3 */
                {8'h31,8'h4b,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SAR,A,4 */
                {8'h31,8'h5b,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SAR,A,5 */
                {8'h31,8'h6b,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SAR,A,6 */
                {8'h31,8'h7b,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SAR,A,7 */
                {8'h31,8'h0f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SARW,AX,0 */
                {8'h31,8'h1f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SARW,AX,1 */
                {8'h31,8'h2f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SARW,AX,2 */
                {8'h31,8'h3f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SARW,AX,3 */
                {8'h31,8'h4f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SARW,AX,4 */
                {8'h31,8'h5f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SARW,AX,5 */
                {8'h31,8'h6f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SARW,AX,6 */
                {8'h31,8'h7f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SARW,AX,7 */
                {8'h31,8'h8f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SARW,AX,8 */
                {8'h31,8'h9f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SARW,AX,9 */
                {8'h31,8'haf,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SARW,AX,10 */
                {8'h31,8'hbf,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SARW,AX,11 */
                {8'h31,8'hcf,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SARW,AX,12 */
                {8'h31,8'hdf,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SARW,AX,13 */
                {8'h31,8'hef,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SARW,AX,14 */
                {8'h31,8'hff,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SARW,AX,15 */
                {8'h61,8'hdb,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ROR,A,1 */
                {8'h61,8'heb,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ROL,A,1 */
                {8'h61,8'hfb,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* RORC,A,1 */
                {8'h61,8'hdc,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ROLC,A,1 */
                {8'h61,8'hee,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ROLWC,AX,1 */
                {8'h61,8'hfe,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ROLWC,BC,1 */
                {8'h71,8'h04,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,saddr.0 */
                {8'h71,8'h14,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,saddr.1 */
                {8'h71,8'h24,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,saddr.2 */
                {8'h71,8'h34,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,saddr.3 */
                {8'h71,8'h44,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,saddr.4 */
                {8'h71,8'h54,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,saddr.5 */
                {8'h71,8'h64,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,saddr.6 */
                {8'h71,8'h74,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,saddr.7 */
                {8'h71,8'h0c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,sfr.0 */
                {8'h71,8'h1c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,sfr.1 */
                {8'h71,8'h2c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,sfr.2 */
                {8'h71,8'h3c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,sfr.3 */
                {8'h71,8'h4c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,sfr.4 */
                {8'h71,8'h5c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,sfr.5 */
                {8'h71,8'h6c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,sfr.6 */
                {8'h71,8'h7c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,sfr.7 */
                {8'h71,8'h8c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,A.0 */
                {8'h71,8'h9c,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,A.1 */
                {8'h71,8'hac,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,A.2 */
                {8'h71,8'hbc,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,A.3 */
                {8'h71,8'hcc,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,A.4 */
                {8'h71,8'hdc,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,A.5 */
                {8'h71,8'hec,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,A.6 */
                {8'h71,8'hfc,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,A.7 */
                {8'h71,8'h84,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,[HL].0 */
                {8'h71,8'h94,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,[HL].1 */
                {8'h71,8'ha4,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,[HL].2 */
                {8'h71,8'hb4,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,[HL].3 */
                {8'h71,8'hc4,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,[HL].4 */
                {8'h71,8'hd4,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,[HL].5 */
                {8'h71,8'he4,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,[HL].6 */
                {8'h71,8'hf4,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* MOV1,CY,[HL].7 */
                {8'h71,8'h05,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,saddr.0 */
                {8'h71,8'h15,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,saddr.1 */
                {8'h71,8'h25,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,saddr.2 */
                {8'h71,8'h35,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,saddr.3 */
                {8'h71,8'h45,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,saddr.4 */
                {8'h71,8'h55,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,saddr.5 */
                {8'h71,8'h65,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,saddr.6 */
                {8'h71,8'h75,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,saddr.7 */
                {8'h71,8'h0d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,sfr.0 */
                {8'h71,8'h1d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,sfr.1 */
                {8'h71,8'h2d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,sfr.2 */
                {8'h71,8'h3d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,sfr.3 */
                {8'h71,8'h4d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,sfr.4 */
                {8'h71,8'h5d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,sfr.5 */
                {8'h71,8'h6d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,sfr.6 */
                {8'h71,8'h7d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,sfr.7 */
                {8'h71,8'h8d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,A.0 */
                {8'h71,8'h9d,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,A.1 */
                {8'h71,8'had,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,A.2 */
                {8'h71,8'hbd,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,A.3 */
                {8'h71,8'hcd,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,A.4 */
                {8'h71,8'hdd,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,A.5 */
                {8'h71,8'hed,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,A.6 */
                {8'h71,8'hfd,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,A.7 */
                {8'h71,8'h85,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,[HL].0 */
                {8'h71,8'h95,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,[HL].1 */
                {8'h71,8'ha5,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,[HL].2 */
                {8'h71,8'hb5,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,[HL].3 */
                {8'h71,8'hc5,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,[HL].4 */
                {8'h71,8'hd5,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,[HL].5 */
                {8'h71,8'he5,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,[HL].6 */
                {8'h71,8'hf5,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* AND1,CY,[HL].7 */
                {8'h71,8'h06,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,saddr.0 */
                {8'h71,8'h16,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,saddr.1 */
                {8'h71,8'h26,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,saddr.2 */
                {8'h71,8'h36,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,saddr.3 */
                {8'h71,8'h46,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,saddr.4 */
                {8'h71,8'h56,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,saddr.5 */
                {8'h71,8'h66,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,saddr.6 */
                {8'h71,8'h76,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,saddr.7 */
                {8'h71,8'h0e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,sfr.0 */
                {8'h71,8'h1e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,sfr.1 */
                {8'h71,8'h2e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,sfr.2 */
                {8'h71,8'h3e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,sfr.3 */
                {8'h71,8'h4e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,sfr.4 */
                {8'h71,8'h5e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,sfr.5 */
                {8'h71,8'h6e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,sfr.6 */
                {8'h71,8'h7e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,sfr.7 */
                {8'h71,8'h8e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,A.0 */
                {8'h71,8'h9e,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,A.1 */
                {8'h71,8'hae,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,A.2 */
                {8'h71,8'hbe,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,A.3 */
                {8'h71,8'hce,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,A.4 */
                {8'h71,8'hde,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,A.5 */
                {8'h71,8'hee,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,A.6 */
                {8'h71,8'hfe,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,A.7 */
                {8'h71,8'h86,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,[HL].0 */
                {8'h71,8'h96,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,[HL].1 */
                {8'h71,8'ha6,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,[HL].2 */
                {8'h71,8'hb6,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,[HL].3 */
                {8'h71,8'hc6,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,[HL].4 */
                {8'h71,8'hd6,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,[HL].5 */
                {8'h71,8'he6,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,[HL].6 */
                {8'h71,8'hf6,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* OR1,CY,[HL].7 */
                {8'h71,8'h07,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,saddr.0 */
                {8'h71,8'h17,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,saddr.1 */
                {8'h71,8'h27,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,saddr.2 */
                {8'h71,8'h37,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,saddr.3 */
                {8'h71,8'h47,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,saddr.4 */
                {8'h71,8'h57,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,saddr.5 */
                {8'h71,8'h67,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,saddr.6 */
                {8'h71,8'h77,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,saddr.7 */
                {8'h71,8'h0f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,sfr.0 */
                {8'h71,8'h1f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,sfr.1 */
                {8'h71,8'h2f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,sfr.2 */
                {8'h71,8'h3f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,sfr.3 */
                {8'h71,8'h4f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,sfr.4 */
                {8'h71,8'h5f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,sfr.5 */
                {8'h71,8'h6f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,sfr.6 */
                {8'h71,8'h7f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,sfr.7 */
                {8'h71,8'h8f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,A.0 */
                {8'h71,8'h9f,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,A.1 */
                {8'h71,8'haf,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,A.2 */
                {8'h71,8'hbf,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,A.3 */
                {8'h71,8'hcf,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,A.4 */
                {8'h71,8'hdf,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,A.5 */
                {8'h71,8'hef,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,A.6 */
                {8'h71,8'hff,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,A.7 */
                {8'h71,8'h87,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,[HL].0 */
                {8'h71,8'h97,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,[HL].1 */
                {8'h71,8'ha7,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,[HL].2 */
                {8'h71,8'hb7,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,[HL].3 */
                {8'h71,8'hc7,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,[HL].4 */
                {8'h71,8'hd7,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,[HL].5 */
                {8'h71,8'he7,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,[HL].6 */
                {8'h71,8'hf7,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* XOR1,CY,[HL].7 */
                {8'h71,8'h80,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SET1,,CY */
                {8'h71,8'h88,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CLR1,,CY */
                {8'h71,8'hc0,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* NOT1,,CY */
                {8'h61,8'hec,2'b01} : dec_CY_enable_adrstage = 1'b1;  /* RETB,, */
                {8'h61,8'hfc,2'b01} : dec_CY_enable_adrstage = 1'b1;  /* RETI,, */
                {8'h61,8'hcd,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* POP,,PSW */
                {8'h61,8'h19,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,A,A */
                {8'h61,8'h39,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,A,A */
                {8'h61,8'h83,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADD,A,[HL+C] */
                {8'h61,8'h93,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* ADDC,A,[HL+C] */
                {8'h61,8'ha3,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUB,A,[HL+C] */
                {8'h61,8'hb3,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SUBC,A,[HL+C] */
                {8'h71,8'h90,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SET1,,CY */
                {8'h71,8'ha0,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SET1,,CY */
                {8'h71,8'hb0,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SET1,,CY */
                {8'h71,8'hd0,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* NOT1,,CY */
                {8'h71,8'he0,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* NOT1,,CY */
                {8'h71,8'hf0,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* NOT1,,CY */
                {8'h71,8'h98,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CLR1,,CY */
                {8'h71,8'ha8,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CLR1,,CY */
                {8'h71,8'hb8,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* CLR1,,CY */
                {8'h71,8'hc8,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* NOT1,,CY */
                {8'h71,8'hd8,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* NOT1,,CY */
                {8'h71,8'he8,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* NOT1,,CY */
                {8'h71,8'hf8,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* NOT1,,CY */
                {8'h31,8'h8a,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHR,A,0 */
                {8'h31,8'h9a,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHR,A,1 */
                {8'h31,8'haa,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHR,A,2 */
                {8'h31,8'hba,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHR,A,3 */
                {8'h31,8'hca,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHR,A,4 */
                {8'h31,8'hda,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHR,A,5 */
                {8'h31,8'hea,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHR,A,6 */
                {8'h31,8'hfa,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHR,A,7 */
                {8'h31,8'h89,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,A,0 */
                {8'h31,8'h99,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,A,1 */
                {8'h31,8'ha9,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,A,2 */
                {8'h31,8'hb9,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,A,3 */
                {8'h31,8'hc9,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,A,4 */
                {8'h31,8'hd9,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,A,5 */
                {8'h31,8'he9,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,A,6 */
                {8'h31,8'hf9,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,A,7 */
                {8'h31,8'h88,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,B,0 */
                {8'h31,8'h98,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,B,1 */
                {8'h31,8'ha8,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,B,2 */
                {8'h31,8'hb8,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,B,3 */
                {8'h31,8'hc8,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,B,4 */
                {8'h31,8'hd8,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,B,5 */
                {8'h31,8'he8,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,B,6 */
                {8'h31,8'hf8,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,B,7 */
                {8'h31,8'h87,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,C,0 */
                {8'h31,8'h97,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,C,1 */
                {8'h31,8'ha7,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,C,2 */
                {8'h31,8'hb7,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,C,3 */
                {8'h31,8'hc7,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,C,4 */
                {8'h31,8'hd7,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,C,5 */
                {8'h31,8'he7,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,C,6 */
                {8'h31,8'hf7,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SHL,C,7 */
                {8'h31,8'h8b,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SAR,A,0 */
                {8'h31,8'h9b,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SAR,A,1 */
                {8'h31,8'hab,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SAR,A,2 */
                {8'h31,8'hbb,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SAR,A,3 */
                {8'h31,8'hcb,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SAR,A,4 */
                {8'h31,8'hdb,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SAR,A,5 */
                {8'h31,8'heb,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SAR,A,6 */
                {8'h31,8'hfb,2'bxx} : dec_CY_enable_adrstage = 1'b1;  /* SAR,A,7 */
                default : dec_CY_enable_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_CY_enable <= 1'b0;
        else if(cpuen) dec_CY_enable <= dec_CY_enable_adrstage;
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*����ADD,ADDC,SUB,SUBC,INC,DEC��						*/
/*���������������ꥢ�������黻�򣲥���å��ܤ��飱����å��ܤ��ѹ�		*/
/*------------------------------------------------------------------------------*/

    output dec_AC_enable;
    reg    dec_AC_enable, dec_AC_enable_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1|| skpack == 1'b1) begin
            dec_AC_enable_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h0c,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,A,#byte */
                {8'h0a,8'hxx,2'bx0} : dec_AC_enable_adrstage = 1'b1;  /* ADD,saddr,#byte */
                {8'h61,8'h08,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,A,X */
                {8'h61,8'h0a,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,A,C */
                {8'h61,8'h0b,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,A,B */
                {8'h61,8'h0c,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,A,E */
                {8'h61,8'h0d,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,A,D */
                {8'h61,8'h0e,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,A,L */
                {8'h61,8'h0f,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,A,H */
                {8'h61,8'h00,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,X,A */
                {8'h61,8'h01,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,A,A */
                {8'h61,8'h02,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,C,A */
                {8'h61,8'h03,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,B,A */
                {8'h61,8'h04,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,E,A */
                {8'h61,8'h05,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,D,A */
                {8'h61,8'h06,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,L,A */
                {8'h61,8'h07,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,H,A */
                {8'h0b,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,A,saddr */
                {8'h0f,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,A,!addr16 */
                {8'h0d,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,A,[HL] */
                {8'h0e,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,A,[HL+byte] */
                {8'h61,8'h80,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,A,[HL+B] */
                {8'h61,8'h82,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,A,[HL+C] */
                {8'h1c,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,A,#byte */
                {8'h1a,8'hxx,2'bx0} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,saddr,#byte */
                {8'h61,8'h18,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,A,X */
                {8'h61,8'h1a,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,A,C */
                {8'h61,8'h1b,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,A,B */
                {8'h61,8'h1c,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,A,E */
                {8'h61,8'h1d,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,A,D */
                {8'h61,8'h1e,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,A,L */
                {8'h61,8'h1f,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,A,H */
                {8'h61,8'h10,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,X,A */
                {8'h61,8'h11,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,A,A */
                {8'h61,8'h12,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,C,A */
                {8'h61,8'h13,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,B,A */
                {8'h61,8'h14,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,E,A */
                {8'h61,8'h15,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,D,A */
                {8'h61,8'h16,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,L,A */
                {8'h61,8'h17,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,H,A */
                {8'h1b,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,A,saddr */
                {8'h1f,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,A,!addr16 */
                {8'h1d,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,A,[HL] */
                {8'h1e,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,A,[HL+byte] */
                {8'h61,8'h90,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,A,[HL+B] */
                {8'h61,8'h92,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,A,[HL+C] */
                {8'h2c,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,A,#byte */
                {8'h2a,8'hxx,2'bx0} : dec_AC_enable_adrstage = 1'b1;  /* SUB,saddr,#byte */
                {8'h61,8'h28,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,A,X */
                {8'h61,8'h2a,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,A,C */
                {8'h61,8'h2b,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,A,B */
                {8'h61,8'h2c,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,A,E */
                {8'h61,8'h2d,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,A,D */
                {8'h61,8'h2e,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,A,L */
                {8'h61,8'h2f,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,A,H */
                {8'h61,8'h20,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,X,A */
                {8'h61,8'h21,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,A,A */
                {8'h61,8'h22,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,C,A */
                {8'h61,8'h23,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,B,A */
                {8'h61,8'h24,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,E,A */
                {8'h61,8'h25,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,D,A */
                {8'h61,8'h26,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,L,A */
                {8'h61,8'h27,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,H,A */
                {8'h2b,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,A,saddr */
                {8'h2f,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,A,!addr16 */
                {8'h2d,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,A,[HL] */
                {8'h2e,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,A,[HL+byte] */
                {8'h61,8'ha0,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,A,[HL+B] */
                {8'h61,8'ha2,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,A,[HL+C] */
                {8'h3c,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,A,#byte */
                {8'h3a,8'hxx,2'bx0} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,saddr,#byte */
                {8'h61,8'h38,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,A,X */
                {8'h61,8'h3a,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,A,C */
                {8'h61,8'h3b,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,A,B */
                {8'h61,8'h3c,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,A,E */
                {8'h61,8'h3d,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,A,D */
                {8'h61,8'h3e,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,A,L */
                {8'h61,8'h3f,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,A,H */
                {8'h61,8'h30,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,X,A */
                {8'h61,8'h31,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,A,A */
                {8'h61,8'h32,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,C,A */
                {8'h61,8'h33,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,B,A */
                {8'h61,8'h34,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,E,A */
                {8'h61,8'h35,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,D,A */
                {8'h61,8'h36,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,L,A */
                {8'h61,8'h37,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,H,A */
                {8'h3b,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,A,saddr */
                {8'h3f,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,A,!addr16 */
                {8'h3d,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,A,[HL] */
                {8'h3e,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,A,[HL+byte] */
                {8'h61,8'hb0,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,A,[HL+B] */
                {8'h61,8'hb2,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,A,[HL+C] */
                {8'h4c,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,A,#byte */
                {8'h4a,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,saddr,#byte */
                {8'h40,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,!addr16,#byte */
                {8'h61,8'h48,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,A,X */
                {8'h61,8'h4a,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,A,C */
                {8'h61,8'h4b,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,A,B */
                {8'h61,8'h4c,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,A,E */
                {8'h61,8'h4d,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,A,D */
                {8'h61,8'h4e,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,A,L */
                {8'h61,8'h4f,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,A,H */
                {8'h61,8'h40,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,X,A */
                {8'h61,8'h41,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,A,A */
                {8'h61,8'h42,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,C,A */
                {8'h61,8'h43,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,B,A */
                {8'h61,8'h44,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,E,A */
                {8'h61,8'h45,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,D,A */
                {8'h61,8'h46,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,L,A */
                {8'h61,8'h47,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,H,A */
                {8'h4b,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,A,saddr */
                {8'h4f,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,A,!addr16 */
                {8'h4d,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,A,[HL] */
                {8'h4e,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,A,[HL+byte] */
                {8'h61,8'hc0,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,A,[HL+B] */
                {8'h61,8'hc2,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP,A,[HL+C] */
                {8'h61,8'hde,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMPS,X,[HL+byte] */
                {8'hd1,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP0,,A */
                {8'hd0,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP0,,X */
                {8'hd3,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP0,,B */
                {8'hd2,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP0,,C */
                {8'hd4,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP0,,saddr */
                {8'hd5,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMP0,,!addr16 */
                {8'h04,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDW,AX,#word */
                {8'h01,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDW,AX,AX */
                {8'h03,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDW,AX,BC */
                {8'h05,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDW,AX,DE */
                {8'h07,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDW,AX,HL */
                {8'h06,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDW,AX,saddrp */
                {8'h02,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDW,AX,!addr16 */
                {8'h61,8'h09,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDW,AX,[HL+byte] */
                {8'h24,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBW,AX,#word */
                {8'h21,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBW,AX,AX */
                {8'h23,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBW,AX,BC */
                {8'h25,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBW,AX,DE */
                {8'h27,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBW,AX,HL */
                {8'h26,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBW,AX,saddrp */
                {8'h22,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBW,AX,!addr16 */
                {8'h61,8'h29,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBW,AX,[HL+byte] */
                {8'h44,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMPW,AX,#word */
                {8'h43,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMPW,AX,BC */
                {8'h45,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMPW,AX,DE */
                {8'h47,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMPW,AX,HL */
                {8'h46,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMPW,AX,saddrp */
                {8'h42,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMPW,AX,!addr16 */
                {8'h61,8'h49,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* CMPW,AX,[HL+byte] */
                {8'h80,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* INC,,X */
                {8'h81,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* INC,,A */
                {8'h82,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* INC,,C */
                {8'h83,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* INC,,B */
                {8'h84,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* INC,,E */
                {8'h85,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* INC,,D */
                {8'h86,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* INC,,L */
                {8'h87,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* INC,,H */
                {8'ha4,8'hxx,2'bx0} : dec_AC_enable_adrstage = 1'b1;  /* INC,,saddr */
                {8'ha0,8'hxx,2'bx0} : dec_AC_enable_adrstage = 1'b1;  /* INC,,!addr16 */
                {8'h61,8'h59,2'bx0} : dec_AC_enable_adrstage = 1'b1;  /* INC,,[HL+byte] */
                {8'h90,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* DEC,,X */
                {8'h91,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* DEC,,A */
                {8'h92,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* DEC,,C */
                {8'h93,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* DEC,,B */
                {8'h94,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* DEC,,E */
                {8'h95,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* DEC,,D */
                {8'h96,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* DEC,,L */
                {8'h97,8'hxx,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* DEC,,H */
                {8'hb4,8'hxx,2'bx0} : dec_AC_enable_adrstage = 1'b1;  /* DEC,,saddr */
                {8'hb0,8'hxx,2'bx0} : dec_AC_enable_adrstage = 1'b1;  /* DEC,,!addr16 */
                {8'h61,8'h69,2'bx0} : dec_AC_enable_adrstage = 1'b1;  /* DEC,,[HL+byte] */
                {8'h61,8'hec,2'b01} : dec_AC_enable_adrstage = 1'b1;  /* RETB,, */
                {8'h61,8'hfc,2'b01} : dec_AC_enable_adrstage = 1'b1;  /* RETI,, */
                {8'h61,8'hcd,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* POP,,PSW */
                {8'h61,8'h19,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,A,A */
                {8'h61,8'h39,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,A,A */
                {8'h61,8'h83,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADD,A,[HL+C] */
                {8'h61,8'h93,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* ADDC,A,[HL+C] */
                {8'h61,8'ha3,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUB,A,[HL+C] */
                {8'h61,8'hb3,2'bxx} : dec_AC_enable_adrstage = 1'b1;  /* SUBC,A,[HL+C] */
                default : dec_AC_enable_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_AC_enable <= 1'b0;
        else if(cpuen) dec_AC_enable <= dec_AC_enable_adrstage;
    end
    output dec_IE_enable;
    reg    dec_IE_enable, dec_IE_enable_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1) begin
            dec_IE_enable_adrstage = 1'b0;
        end else if(ivack == 1'b1) begin
            casex ({stage_adr})  
                {2'b10} : dec_IE_enable_adrstage = 1'b1;  /* Interrupt */
                default : dec_IE_enable_adrstage = 1'b0;
            endcase
        end else if(skpack == 1'b1) begin
            dec_IE_enable_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hec,2'b01} : dec_IE_enable_adrstage = 1'b1;  /* RETB,, */
                {8'h61,8'hfc,2'b01} : dec_IE_enable_adrstage = 1'b1;  /* RETI,, */
                {8'h61,8'hcd,2'bxx} : dec_IE_enable_adrstage = 1'b1;  /* POP,,PSW */
                default : dec_IE_enable_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_IE_enable <= 1'b0;
        else if(cpuen) dec_IE_enable <= dec_IE_enable_adrstage;
    end
    output dec_ISP_enable;
    reg    dec_ISP_enable, dec_ISP_enable_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1|| skpack == 1'b1) begin
            dec_ISP_enable_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hec,2'b01} : dec_ISP_enable_adrstage = 1'b1;  /* RETB,, */
                {8'h61,8'hfc,2'b01} : dec_ISP_enable_adrstage = 1'b1;  /* RETI,, */
                {8'h61,8'hcd,2'bxx} : dec_ISP_enable_adrstage = 1'b1;  /* POP,,PSW */
                default : dec_ISP_enable_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_ISP_enable <= 1'b0;
        else if(cpuen) dec_ISP_enable <= dec_ISP_enable_adrstage;
    end
    output dec_RBS_enable;
    reg    dec_RBS_enable, dec_RBS_enable_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1|| skpack == 1'b1) begin
            dec_RBS_enable_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hec,2'b01} : dec_RBS_enable_adrstage = 1'b1;  /* RETB,, */
                {8'h61,8'hfc,2'b01} : dec_RBS_enable_adrstage = 1'b1;  /* RETI,, */
                {8'h61,8'hcd,2'bxx} : dec_RBS_enable_adrstage = 1'b1;  /* POP,,PSW */
                {8'h61,8'hcf,2'bxx} : dec_RBS_enable_adrstage = 1'b1;  /* SEL,,RB0 */
                {8'h61,8'hdf,2'bxx} : dec_RBS_enable_adrstage = 1'b1;  /* SEL,,RB1 */
                {8'h61,8'hef,2'bxx} : dec_RBS_enable_adrstage = 1'b1;  /* SEL,,RB2 */
                {8'h61,8'hff,2'bxx} : dec_RBS_enable_adrstage = 1'b1;  /* SEL,,RB3 */
                default : dec_RBS_enable_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_RBS_enable <= 1'b0;
        else if(cpuen) dec_RBS_enable <= dec_RBS_enable_adrstage;
    end
    output dec_NMIS_enable;
    reg    dec_NMIS_enable, dec_NMIS_enable_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1|| skpack == 1'b1) begin
            dec_NMIS_enable_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hfc,2'b01} : dec_NMIS_enable_adrstage = 1'b1;  /* RETI,, */
                default : dec_NMIS_enable_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_NMIS_enable <= 1'b0;
        else if(cpuen) dec_NMIS_enable <= dec_NMIS_enable_adrstage;
    end
    output dec_buf0_enable;
    reg    dec_buf0_enable, dec_buf0_enable_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1|| skpack == 1'b1) begin
            dec_buf0_enable_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'ha8,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* XCH,A,saddr */
                {8'h61,8'hab,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* XCH,A,sfr */
                {8'h61,8'haa,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* XCH,A,!addr16 */
                {8'h61,8'hae,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* XCH,A,[DE] */
                {8'h61,8'haf,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* XCH,A,[DE+byte] */
                {8'h61,8'hac,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* XCH,A,[HL] */
                {8'h61,8'had,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* XCH,A,[HL+byte] */
                {8'h61,8'hb9,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* XCH,A,[HL+B] */
                {8'h61,8'ha9,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* XCH,A,[HL+C] */
                {8'h0a,8'hxx,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* ADD,saddr,#byte */
                {8'h1a,8'hxx,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* ADDC,saddr,#byte */
                {8'h2a,8'hxx,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SUB,saddr,#byte */
                {8'h3a,8'hxx,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SUBC,saddr,#byte */
                {8'h5a,8'hxx,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* AND,saddr,#byte */
                {8'h6a,8'hxx,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* OR,saddr,#byte */
                {8'h7a,8'hxx,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* XOR,saddr,#byte */
                {8'ha4,8'hxx,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* INC,,saddr */
                {8'ha0,8'hxx,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* INC,,!addr16 */
                {8'h61,8'h59,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* INC,,[HL+byte] */
                {8'hb4,8'hxx,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* DEC,,saddr */
                {8'hb0,8'hxx,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* DEC,,!addr16 */
                {8'h61,8'h69,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* DEC,,[HL+byte] */
                {8'ha6,8'hxx,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* INCW,,saddrp */
                {8'ha2,8'hxx,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* INCW,,!addr16 */
                {8'h61,8'h79,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* INCW,,[HL+byte] */
                {8'hb6,8'hxx,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* DECW,,saddrp */
                {8'hb2,8'hxx,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* DECW,,!addr16 */
                {8'h61,8'h89,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* DECW,,[HL+byte] */
                {8'h71,8'h01,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,saddr.0,CY */
                {8'h71,8'h11,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,saddr.1,CY */
                {8'h71,8'h21,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,saddr.2,CY */
                {8'h71,8'h31,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,saddr.3,CY */
                {8'h71,8'h41,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,saddr.4,CY */
                {8'h71,8'h51,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,saddr.5,CY */
                {8'h71,8'h61,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,saddr.6,CY */
                {8'h71,8'h71,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,saddr.7,CY */
                {8'h71,8'h09,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,sfr.0,CY */
                {8'h71,8'h19,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,sfr.1,CY */
                {8'h71,8'h29,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,sfr.2,CY */
                {8'h71,8'h39,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,sfr.3,CY */
                {8'h71,8'h49,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,sfr.4,CY */
                {8'h71,8'h59,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,sfr.5,CY */
                {8'h71,8'h69,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,sfr.6,CY */
                {8'h71,8'h79,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,sfr.7,CY */
                {8'h71,8'h81,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,[HL].0,CY */
                {8'h71,8'h91,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,[HL].1,CY */
                {8'h71,8'ha1,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,[HL].2,CY */
                {8'h71,8'hb1,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,[HL].3,CY */
                {8'h71,8'hc1,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,[HL].4,CY */
                {8'h71,8'hd1,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,[HL].5,CY */
                {8'h71,8'he1,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,[HL].6,CY */
                {8'h71,8'hf1,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* MOV1,[HL].7,CY */
                {8'h71,8'h02,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,saddr.0 */
                {8'h71,8'h12,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,saddr.1 */
                {8'h71,8'h22,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,saddr.2 */
                {8'h71,8'h32,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,saddr.3 */
                {8'h71,8'h42,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,saddr.4 */
                {8'h71,8'h52,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,saddr.5 */
                {8'h71,8'h62,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,saddr.6 */
                {8'h71,8'h72,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,saddr.7 */
                {8'h71,8'h0a,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,sfr.0 */
                {8'h71,8'h1a,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,sfr.1 */
                {8'h71,8'h2a,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,sfr.2 */
                {8'h71,8'h3a,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,sfr.3 */
                {8'h71,8'h4a,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,sfr.4 */
                {8'h71,8'h5a,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,sfr.5 */
                {8'h71,8'h6a,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,sfr.6 */
                {8'h71,8'h7a,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,sfr.7 */
                {8'h71,8'h00,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,!addr16.0 */
                {8'h71,8'h10,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,!addr16.1 */
                {8'h71,8'h20,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,!addr16.2 */
                {8'h71,8'h30,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,!addr16.3 */
                {8'h71,8'h40,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,!addr16.4 */
                {8'h71,8'h50,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,!addr16.5 */
                {8'h71,8'h60,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,!addr16.6 */
                {8'h71,8'h70,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,!addr16.7 */
                {8'h71,8'h82,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,[HL].0 */
                {8'h71,8'h92,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,[HL].1 */
                {8'h71,8'ha2,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,[HL].2 */
                {8'h71,8'hb2,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,[HL].3 */
                {8'h71,8'hc2,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,[HL].4 */
                {8'h71,8'hd2,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,[HL].5 */
                {8'h71,8'he2,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,[HL].6 */
                {8'h71,8'hf2,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* SET1,,[HL].7 */
                {8'h71,8'h03,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,saddr.0 */
                {8'h71,8'h13,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,saddr.1 */
                {8'h71,8'h23,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,saddr.2 */
                {8'h71,8'h33,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,saddr.3 */
                {8'h71,8'h43,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,saddr.4 */
                {8'h71,8'h53,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,saddr.5 */
                {8'h71,8'h63,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,saddr.6 */
                {8'h71,8'h73,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,saddr.7 */
                {8'h71,8'h0b,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,sfr.0 */
                {8'h71,8'h1b,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,sfr.1 */
                {8'h71,8'h2b,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,sfr.2 */
                {8'h71,8'h3b,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,sfr.3 */
                {8'h71,8'h4b,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,sfr.4 */
                {8'h71,8'h5b,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,sfr.5 */
                {8'h71,8'h6b,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,sfr.6 */
                {8'h71,8'h7b,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,sfr.7 */
                {8'h71,8'h08,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,!addr16.0 */
                {8'h71,8'h18,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,!addr16.1 */
                {8'h71,8'h28,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,!addr16.2 */
                {8'h71,8'h38,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,!addr16.3 */
                {8'h71,8'h48,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,!addr16.4 */
                {8'h71,8'h58,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,!addr16.5 */
                {8'h71,8'h68,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,!addr16.6 */
                {8'h71,8'h78,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,!addr16.7 */
                {8'h71,8'h83,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,[HL].0 */
                {8'h71,8'h93,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,[HL].1 */
                {8'h71,8'ha3,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,[HL].2 */
                {8'h71,8'hb3,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,[HL].3 */
                {8'h71,8'hc3,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,[HL].4 */
                {8'h71,8'hd3,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,[HL].5 */
                {8'h71,8'he3,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,[HL].6 */
                {8'h71,8'hf3,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* CLR1,,[HL].7 */
                {8'hd7,8'hxx,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* RET,, */
                {8'h61,8'hec,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* RETB,, */
                {8'h61,8'hfc,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* RETI,, */
                {8'h31,8'h02,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,saddr.0,$addr8 */
                {8'h31,8'h12,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,saddr.1,$addr8 */
                {8'h31,8'h22,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,saddr.2,$addr8 */
                {8'h31,8'h32,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,saddr.3,$addr8 */
                {8'h31,8'h42,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,saddr.4,$addr8 */
                {8'h31,8'h52,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,saddr.5,$addr8 */
                {8'h31,8'h62,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,saddr.6,$addr8 */
                {8'h31,8'h72,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,saddr.7,$addr8 */
                {8'h31,8'h82,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,sfr.0,$addr8 */
                {8'h31,8'h92,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,sfr.1,$addr8 */
                {8'h31,8'ha2,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,sfr.2,$addr8 */
                {8'h31,8'hb2,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,sfr.3,$addr8 */
                {8'h31,8'hc2,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,sfr.4,$addr8 */
                {8'h31,8'hd2,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,sfr.5,$addr8 */
                {8'h31,8'he2,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,sfr.6,$addr8 */
                {8'h31,8'hf2,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,sfr.7,$addr8 */
                {8'h31,8'h03,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,A.0,$addr8 */
                {8'h31,8'h13,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,A.1,$addr8 */
                {8'h31,8'h23,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,A.2,$addr8 */
                {8'h31,8'h33,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,A.3,$addr8 */
                {8'h31,8'h43,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,A.4,$addr8 */
                {8'h31,8'h53,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,A.5,$addr8 */
                {8'h31,8'h63,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,A.6,$addr8 */
                {8'h31,8'h73,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,A.7,$addr8 */
                {8'h31,8'h83,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,[HL].0,$addr8 */
                {8'h31,8'h93,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,[HL].1,$addr8 */
                {8'h31,8'ha3,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,[HL].2,$addr8 */
                {8'h31,8'hb3,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,[HL].3,$addr8 */
                {8'h31,8'hc3,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,[HL].4,$addr8 */
                {8'h31,8'hd3,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,[HL].5,$addr8 */
                {8'h31,8'he3,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,[HL].6,$addr8 */
                {8'h31,8'hf3,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BT,[HL].7,$addr8 */
                {8'h31,8'h04,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,saddr.0,$addr8 */
                {8'h31,8'h14,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,saddr.1,$addr8 */
                {8'h31,8'h24,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,saddr.2,$addr8 */
                {8'h31,8'h34,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,saddr.3,$addr8 */
                {8'h31,8'h44,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,saddr.4,$addr8 */
                {8'h31,8'h54,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,saddr.5,$addr8 */
                {8'h31,8'h64,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,saddr.6,$addr8 */
                {8'h31,8'h74,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,saddr.7,$addr8 */
                {8'h31,8'h84,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,sfr.0,$addr8 */
                {8'h31,8'h94,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,sfr.1,$addr8 */
                {8'h31,8'ha4,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,sfr.2,$addr8 */
                {8'h31,8'hb4,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,sfr.3,$addr8 */
                {8'h31,8'hc4,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,sfr.4,$addr8 */
                {8'h31,8'hd4,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,sfr.5,$addr8 */
                {8'h31,8'he4,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,sfr.6,$addr8 */
                {8'h31,8'hf4,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,sfr.7,$addr8 */
                {8'h31,8'h05,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,A.0,$addr8 */
                {8'h31,8'h15,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,A.1,$addr8 */
                {8'h31,8'h25,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,A.2,$addr8 */
                {8'h31,8'h35,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,A.3,$addr8 */
                {8'h31,8'h45,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,A.4,$addr8 */
                {8'h31,8'h55,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,A.5,$addr8 */
                {8'h31,8'h65,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,A.6,$addr8 */
                {8'h31,8'h75,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,A.7,$addr8 */
                {8'h31,8'h85,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,[HL].0,$addr8 */
                {8'h31,8'h95,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,[HL].1,$addr8 */
                {8'h31,8'ha5,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,[HL].2,$addr8 */
                {8'h31,8'hb5,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,[HL].3,$addr8 */
                {8'h31,8'hc5,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,[HL].4,$addr8 */
                {8'h31,8'hd5,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,[HL].5,$addr8 */
                {8'h31,8'he5,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,[HL].6,$addr8 */
                {8'h31,8'hf5,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BF,[HL].7,$addr8 */
                {8'h31,8'h00,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,saddr.0,$addr8 */
                {8'h31,8'h00,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,saddr.0,$addr8 */
                {8'h31,8'h10,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,saddr.1,$addr8 */
                {8'h31,8'h10,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,saddr.1,$addr8 */
                {8'h31,8'h20,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,saddr.2,$addr8 */
                {8'h31,8'h20,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,saddr.2,$addr8 */
                {8'h31,8'h30,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,saddr.3,$addr8 */
                {8'h31,8'h30,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,saddr.3,$addr8 */
                {8'h31,8'h40,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,saddr.4,$addr8 */
                {8'h31,8'h40,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,saddr.4,$addr8 */
                {8'h31,8'h50,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,saddr.5,$addr8 */
                {8'h31,8'h50,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,saddr.5,$addr8 */
                {8'h31,8'h60,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,saddr.6,$addr8 */
                {8'h31,8'h60,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,saddr.6,$addr8 */
                {8'h31,8'h70,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,saddr.7,$addr8 */
                {8'h31,8'h70,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,saddr.7,$addr8 */
                {8'h31,8'h80,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,sfr.0,$addr8 */
                {8'h31,8'h80,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,sfr.0,$addr8 */
                {8'h31,8'h90,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,sfr.1,$addr8 */
                {8'h31,8'h90,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,sfr.1,$addr8 */
                {8'h31,8'ha0,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,sfr.2,$addr8 */
                {8'h31,8'ha0,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,sfr.2,$addr8 */
                {8'h31,8'hb0,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,sfr.3,$addr8 */
                {8'h31,8'hb0,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,sfr.3,$addr8 */
                {8'h31,8'hc0,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,sfr.4,$addr8 */
                {8'h31,8'hc0,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,sfr.4,$addr8 */
                {8'h31,8'hd0,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,sfr.5,$addr8 */
                {8'h31,8'hd0,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,sfr.5,$addr8 */
                {8'h31,8'he0,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,sfr.6,$addr8 */
                {8'h31,8'he0,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,sfr.6,$addr8 */
                {8'h31,8'hf0,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,sfr.7,$addr8 */
                {8'h31,8'hf0,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,sfr.7,$addr8 */
                {8'h31,8'h01,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,A.0,$addr8 */
                {8'h31,8'h11,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,A.1,$addr8 */
                {8'h31,8'h21,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,A.2,$addr8 */
                {8'h31,8'h31,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,A.3,$addr8 */
                {8'h31,8'h41,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,A.4,$addr8 */
                {8'h31,8'h51,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,A.5,$addr8 */
                {8'h31,8'h61,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,A.6,$addr8 */
                {8'h31,8'h71,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,A.7,$addr8 */
                {8'h31,8'h81,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,[HL].0,$addr8 */
                {8'h31,8'h81,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,[HL].0,$addr8 */
                {8'h31,8'h91,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,[HL].1,$addr8 */
                {8'h31,8'h91,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,[HL].1,$addr8 */
                {8'h31,8'ha1,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,[HL].2,$addr8 */
                {8'h31,8'ha1,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,[HL].2,$addr8 */
                {8'h31,8'hb1,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,[HL].3,$addr8 */
                {8'h31,8'hb1,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,[HL].3,$addr8 */
                {8'h31,8'hc1,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,[HL].4,$addr8 */
                {8'h31,8'hc1,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,[HL].4,$addr8 */
                {8'h31,8'hd1,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,[HL].5,$addr8 */
                {8'h31,8'hd1,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,[HL].5,$addr8 */
                {8'h31,8'he1,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,[HL].6,$addr8 */
                {8'h31,8'he1,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,[HL].6,$addr8 */
                {8'h31,8'hf1,2'b00} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,[HL].7,$addr8 */
                {8'h31,8'hf1,2'b01} : dec_buf0_enable_adrstage = 1'b1;  /* BTCLR,[HL].7,$addr8 */
                {8'h61,8'hbb,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* XCH,A,sfr */
                {8'h61,8'hba,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* XCH,A,!addr16 */
                {8'h61,8'hbe,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* XCH,A,[DE] */
                {8'h61,8'hbf,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* XCH,A,[DE+byte] */
                {8'h61,8'hbc,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* XCH,A,[HL] */
                {8'h61,8'hbd,2'bx0} : dec_buf0_enable_adrstage = 1'b1;  /* XCH,A,[HL+byte] */
                default : dec_buf0_enable_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_buf0_enable <= 1'b0;
        else if(cpuen) dec_buf0_enable <= dec_buf0_enable_adrstage;
    end
    output dec_buf1_enable;
    reg    dec_buf1_enable, dec_buf1_enable_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1|| skpack == 1'b1) begin
            dec_buf1_enable_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'ha6,8'hxx,2'bx0} : dec_buf1_enable_adrstage = 1'b1;  /* INCW,,saddrp */
                {8'ha2,8'hxx,2'bx0} : dec_buf1_enable_adrstage = 1'b1;  /* INCW,,!addr16 */
                {8'h61,8'h79,2'bx0} : dec_buf1_enable_adrstage = 1'b1;  /* INCW,,[HL+byte] */
                {8'hb6,8'hxx,2'bx0} : dec_buf1_enable_adrstage = 1'b1;  /* DECW,,saddrp */
                {8'hb2,8'hxx,2'bx0} : dec_buf1_enable_adrstage = 1'b1;  /* DECW,,!addr16 */
                {8'h61,8'h89,2'bx0} : dec_buf1_enable_adrstage = 1'b1;  /* DECW,,[HL+byte] */
                {8'hd7,8'hxx,2'b00} : dec_buf1_enable_adrstage = 1'b1;  /* RET,, */
                {8'h61,8'hec,2'b00} : dec_buf1_enable_adrstage = 1'b1;  /* RETB,, */
                {8'h61,8'hfc,2'b00} : dec_buf1_enable_adrstage = 1'b1;  /* RETI,, */
                default : dec_buf1_enable_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_buf1_enable <= 1'b0;
        else if(cpuen) dec_buf1_enable <= dec_buf1_enable_adrstage;
    end
    output dec_buf2_enable;
    reg    dec_buf2_enable, dec_buf2_enable_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1|| skpack == 1'b1) begin
            dec_buf2_enable_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'hd7,8'hxx,2'b01} : dec_buf2_enable_adrstage = 1'b1;  /* RET,, */
                {8'h61,8'hec,2'b01} : dec_buf2_enable_adrstage = 1'b1;  /* RETB,, */
                {8'h61,8'hfc,2'b01} : dec_buf2_enable_adrstage = 1'b1;  /* RETI,, */
                default : dec_buf2_enable_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_buf2_enable <= 1'b0;
        else if(cpuen) dec_buf2_enable <= dec_buf2_enable_adrstage;
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_cpuwr_enable;
    reg    dec_cpuwr_enable;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(decout_mask == 1'b1) begin
//            dec_cpuwr_enable = 1'b0;
//        end else if(rstvec == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1) begin
            dec_cpuwr_enable = 1'b0;
        end else if(skpack == 1'b1) begin
            dec_cpuwr_enable = 1'b0;
        end else if(ivack == 1'b1) begin
            casex ({stage_adr})  
                {2'b00} : dec_cpuwr_enable = 1'b1;  /* Interrupt */
                {2'b01} : dec_cpuwr_enable = 1'b1;  /* Interrupt */
                default : dec_cpuwr_enable = 1'b0;
            endcase
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'hcd,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOV,saddr,#byte */
                {8'hce,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOV,sfr,#byte */
                {8'hcf,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOV,!addr16,#byte */
                {8'hca,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOV,[DE+byte],#byte */
                {8'hcc,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOV,[HL+byte],#byte */
                {8'h9d,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOV,saddr,A */
                {8'h9e,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOV,sfr,A */
                {8'h9f,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOV,!addr16,A */
                {8'h99,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOV,[DE],A */
                {8'h9a,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOV,[DE+byte],A */
                {8'h9b,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOV,[HL],A */
                {8'h9c,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOV,[HL+byte],A */
                {8'h61,8'hd9,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOV,[HL+B],A */
                {8'h61,8'hf9,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOV,[HL+C],A */
                {8'h19,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOV,word[B],#byte */
                {8'h18,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOV,word[B],A */
                {8'h38,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOV,word[C],#byte */
                {8'h28,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOV,word[C],A */
                {8'h39,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOV,word[BC],#byte */
                {8'h48,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOV,word[BC],A */
                {8'hc8,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOV,[SP+byte],#byte */
                {8'h98,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOV,[SP+byte],A */
                {8'h61,8'hce,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOVS,[HL+byte],X */
                {8'h61,8'ha8,2'bx1} : dec_cpuwr_enable = 1'b1;  /* XCH,A,saddr */
                {8'h61,8'hab,2'bx1} : dec_cpuwr_enable = 1'b1;  /* XCH,A,sfr */
                {8'h61,8'haa,2'bx1} : dec_cpuwr_enable = 1'b1;  /* XCH,A,!addr16 */
                {8'h61,8'hae,2'bx1} : dec_cpuwr_enable = 1'b1;  /* XCH,A,[DE] */
                {8'h61,8'haf,2'bx1} : dec_cpuwr_enable = 1'b1;  /* XCH,A,[DE+byte] */
                {8'h61,8'hac,2'bx1} : dec_cpuwr_enable = 1'b1;  /* XCH,A,[HL] */
                {8'h61,8'had,2'bx1} : dec_cpuwr_enable = 1'b1;  /* XCH,A,[HL+byte] */
                {8'h61,8'hb9,2'bx1} : dec_cpuwr_enable = 1'b1;  /* XCH,A,[HL+B] */
                {8'h61,8'ha9,2'bx1} : dec_cpuwr_enable = 1'b1;  /* XCH,A,[HL+C] */
                {8'he4,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* ONEB,,saddr */
                {8'he5,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* ONEB,,!addr16 */
                {8'hf4,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* CLRB,,saddr */
                {8'hf5,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* CLRB,,!addr16 */
                {8'hc9,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOVW,saddrp,#word */
                {8'hcb,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOVW,sfrp,#word */
                {8'hbd,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOVW,saddrp,AX */
                {8'hbe,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOVW,sfrp,AX */
                {8'hbf,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOVW,!addr16,AX */
                {8'hb9,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOVW,[DE],AX */
                {8'hba,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOVW,[DE+byte],AX */
                {8'hbb,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOVW,[HL],AX */
                {8'hbc,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOVW,[HL+byte],AX */
                {8'h58,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOVW,word[B],AX */
                {8'h68,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOVW,word[C],AX */
                {8'h78,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOVW,word[BC],AX */
                {8'hb8,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* MOVW,[SP+byte],AX */
                {8'h0a,8'hxx,2'bx1} : dec_cpuwr_enable = 1'b1;  /* ADD,saddr,#byte */
                {8'h1a,8'hxx,2'bx1} : dec_cpuwr_enable = 1'b1;  /* ADDC,saddr,#byte */
                {8'h2a,8'hxx,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SUB,saddr,#byte */
                {8'h3a,8'hxx,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SUBC,saddr,#byte */
                {8'h5a,8'hxx,2'bx1} : dec_cpuwr_enable = 1'b1;  /* AND,saddr,#byte */
                {8'h6a,8'hxx,2'bx1} : dec_cpuwr_enable = 1'b1;  /* OR,saddr,#byte */
                {8'h7a,8'hxx,2'bx1} : dec_cpuwr_enable = 1'b1;  /* XOR,saddr,#byte */
                {8'ha4,8'hxx,2'bx1} : dec_cpuwr_enable = 1'b1;  /* INC,,saddr */
                {8'ha0,8'hxx,2'bx1} : dec_cpuwr_enable = 1'b1;  /* INC,,!addr16 */
                {8'h61,8'h59,2'bx1} : dec_cpuwr_enable = 1'b1;  /* INC,,[HL+byte] */
                {8'hb4,8'hxx,2'bx1} : dec_cpuwr_enable = 1'b1;  /* DEC,,saddr */
                {8'hb0,8'hxx,2'bx1} : dec_cpuwr_enable = 1'b1;  /* DEC,,!addr16 */
                {8'h61,8'h69,2'bx1} : dec_cpuwr_enable = 1'b1;  /* DEC,,[HL+byte] */
                {8'ha6,8'hxx,2'bx1} : dec_cpuwr_enable = 1'b1;  /* INCW,,saddrp */
                {8'ha2,8'hxx,2'bx1} : dec_cpuwr_enable = 1'b1;  /* INCW,,!addr16 */
                {8'h61,8'h79,2'bx1} : dec_cpuwr_enable = 1'b1;  /* INCW,,[HL+byte] */
                {8'hb6,8'hxx,2'bx1} : dec_cpuwr_enable = 1'b1;  /* DECW,,saddrp */
                {8'hb2,8'hxx,2'bx1} : dec_cpuwr_enable = 1'b1;  /* DECW,,!addr16 */
                {8'h61,8'h89,2'bx1} : dec_cpuwr_enable = 1'b1;  /* DECW,,[HL+byte] */
                {8'h71,8'h01,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,saddr.0,CY */
                {8'h71,8'h11,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,saddr.1,CY */
                {8'h71,8'h21,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,saddr.2,CY */
                {8'h71,8'h31,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,saddr.3,CY */
                {8'h71,8'h41,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,saddr.4,CY */
                {8'h71,8'h51,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,saddr.5,CY */
                {8'h71,8'h61,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,saddr.6,CY */
                {8'h71,8'h71,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,saddr.7,CY */
                {8'h71,8'h09,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,sfr.0,CY */
                {8'h71,8'h19,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,sfr.1,CY */
                {8'h71,8'h29,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,sfr.2,CY */
                {8'h71,8'h39,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,sfr.3,CY */
                {8'h71,8'h49,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,sfr.4,CY */
                {8'h71,8'h59,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,sfr.5,CY */
                {8'h71,8'h69,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,sfr.6,CY */
                {8'h71,8'h79,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,sfr.7,CY */
                {8'h71,8'h81,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,[HL].0,CY */
                {8'h71,8'h91,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,[HL].1,CY */
                {8'h71,8'ha1,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,[HL].2,CY */
                {8'h71,8'hb1,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,[HL].3,CY */
                {8'h71,8'hc1,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,[HL].4,CY */
                {8'h71,8'hd1,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,[HL].5,CY */
                {8'h71,8'he1,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,[HL].6,CY */
                {8'h71,8'hf1,2'bx1} : dec_cpuwr_enable = 1'b1;  /* MOV1,[HL].7,CY */
                {8'h71,8'h02,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,saddr.0 */
                {8'h71,8'h12,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,saddr.1 */
                {8'h71,8'h22,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,saddr.2 */
                {8'h71,8'h32,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,saddr.3 */
                {8'h71,8'h42,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,saddr.4 */
                {8'h71,8'h52,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,saddr.5 */
                {8'h71,8'h62,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,saddr.6 */
                {8'h71,8'h72,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,saddr.7 */
                {8'h71,8'h0a,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,sfr.0 */
                {8'h71,8'h1a,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,sfr.1 */
                {8'h71,8'h2a,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,sfr.2 */
                {8'h71,8'h3a,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,sfr.3 */
                {8'h71,8'h4a,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,sfr.4 */
                {8'h71,8'h5a,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,sfr.5 */
                {8'h71,8'h6a,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,sfr.6 */
                {8'h71,8'h7a,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,sfr.7 */
                {8'h71,8'h00,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,!addr16.0 */
                {8'h71,8'h10,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,!addr16.1 */
                {8'h71,8'h20,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,!addr16.2 */
                {8'h71,8'h30,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,!addr16.3 */
                {8'h71,8'h40,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,!addr16.4 */
                {8'h71,8'h50,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,!addr16.5 */
                {8'h71,8'h60,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,!addr16.6 */
                {8'h71,8'h70,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,!addr16.7 */
                {8'h71,8'h82,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,[HL].0 */
                {8'h71,8'h92,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,[HL].1 */
                {8'h71,8'ha2,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,[HL].2 */
                {8'h71,8'hb2,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,[HL].3 */
                {8'h71,8'hc2,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,[HL].4 */
                {8'h71,8'hd2,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,[HL].5 */
                {8'h71,8'he2,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,[HL].6 */
                {8'h71,8'hf2,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SET1,,[HL].7 */
                {8'h71,8'h03,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,saddr.0 */
                {8'h71,8'h13,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,saddr.1 */
                {8'h71,8'h23,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,saddr.2 */
                {8'h71,8'h33,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,saddr.3 */
                {8'h71,8'h43,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,saddr.4 */
                {8'h71,8'h53,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,saddr.5 */
                {8'h71,8'h63,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,saddr.6 */
                {8'h71,8'h73,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,saddr.7 */
                {8'h71,8'h0b,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,sfr.0 */
                {8'h71,8'h1b,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,sfr.1 */
                {8'h71,8'h2b,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,sfr.2 */
                {8'h71,8'h3b,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,sfr.3 */
                {8'h71,8'h4b,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,sfr.4 */
                {8'h71,8'h5b,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,sfr.5 */
                {8'h71,8'h6b,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,sfr.6 */
                {8'h71,8'h7b,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,sfr.7 */
                {8'h71,8'h08,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,!addr16.0 */
                {8'h71,8'h18,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,!addr16.1 */
                {8'h71,8'h28,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,!addr16.2 */
                {8'h71,8'h38,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,!addr16.3 */
                {8'h71,8'h48,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,!addr16.4 */
                {8'h71,8'h58,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,!addr16.5 */
                {8'h71,8'h68,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,!addr16.6 */
                {8'h71,8'h78,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,!addr16.7 */
                {8'h71,8'h83,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,[HL].0 */
                {8'h71,8'h93,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,[HL].1 */
                {8'h71,8'ha3,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,[HL].2 */
                {8'h71,8'hb3,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,[HL].3 */
                {8'h71,8'hc3,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,[HL].4 */
                {8'h71,8'hd3,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,[HL].5 */
                {8'h71,8'he3,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,[HL].6 */
                {8'h71,8'hf3,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CLR1,,[HL].7 */
                {8'h61,8'hca,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALL,,AX */
                {8'h61,8'hca,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALL,,AX */
                {8'h61,8'hda,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALL,,BC */
                {8'h61,8'hda,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALL,,BC */
                {8'h61,8'hea,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALL,,DE */
                {8'h61,8'hea,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALL,,DE */
                {8'h61,8'hfa,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALL,,HL */
                {8'h61,8'hfa,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALL,,HL */
                {8'hfe,8'hxx,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALL,,$!addr16 */
                {8'hfe,8'hxx,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALL,,$!addr16 */
                {8'hfd,8'hxx,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALL,,!addr16 */
                {8'hfd,8'hxx,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALL,,!addr16 */
                {8'hfc,8'hxx,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALL,,!!addr20 */
                {8'hfc,8'hxx,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALL,,!!addr20 */
                {8'h61,8'h84,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[0080h] */
                {8'h61,8'h84,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[0080h] */
                {8'h61,8'h94,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[0082h] */
                {8'h61,8'h94,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[0082h] */
                {8'h61,8'ha4,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[0084h] */
                {8'h61,8'ha4,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[0084h] */
                {8'h61,8'hb4,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[0086h] */
                {8'h61,8'hb4,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[0086h] */
                {8'h61,8'hc4,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[0088h] */
                {8'h61,8'hc4,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[0088h] */
                {8'h61,8'hd4,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[008Ah] */
                {8'h61,8'hd4,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[008Ah] */
                {8'h61,8'he4,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[008Ch] */
                {8'h61,8'he4,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[008Ch] */
                {8'h61,8'hf4,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[008Eh] */
                {8'h61,8'hf4,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[008Eh] */
                {8'h61,8'h85,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[0090h] */
                {8'h61,8'h85,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[0090h] */
                {8'h61,8'h95,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[0092h] */
                {8'h61,8'h95,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[0092h] */
                {8'h61,8'ha5,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[0094h] */
                {8'h61,8'ha5,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[0094h] */
                {8'h61,8'hb5,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[0096h] */
                {8'h61,8'hb5,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[0096h] */
                {8'h61,8'hc5,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[0098h] */
                {8'h61,8'hc5,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[0098h] */
                {8'h61,8'hd5,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[009Ah] */
                {8'h61,8'hd5,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[009Ah] */
                {8'h61,8'he5,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[009Ch] */
                {8'h61,8'he5,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[009Ch] */
                {8'h61,8'hf5,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[009Eh] */
                {8'h61,8'hf5,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[009Eh] */
                {8'h61,8'h86,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00A0h] */
                {8'h61,8'h86,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00A0h] */
                {8'h61,8'h96,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00A2h] */
                {8'h61,8'h96,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00A2h] */
                {8'h61,8'ha6,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00A4h] */
                {8'h61,8'ha6,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00A4h] */
                {8'h61,8'hb6,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00A6h] */
                {8'h61,8'hb6,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00A6h] */
                {8'h61,8'hc6,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00A8h] */
                {8'h61,8'hc6,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00A8h] */
                {8'h61,8'hd6,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00AAh] */
                {8'h61,8'hd6,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00AAh] */
                {8'h61,8'he6,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00ACh] */
                {8'h61,8'he6,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00ACh] */
                {8'h61,8'hf6,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00AEh] */
                {8'h61,8'hf6,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00AEh] */
                {8'h61,8'h87,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00B0h] */
                {8'h61,8'h87,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00B0h] */
                {8'h61,8'h97,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00B2h] */
                {8'h61,8'h97,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00B2h] */
                {8'h61,8'ha7,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00B4h] */
                {8'h61,8'ha7,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00B4h] */
                {8'h61,8'hb7,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00B6h] */
                {8'h61,8'hb7,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00B6h] */
                {8'h61,8'hc7,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00B8h] */
                {8'h61,8'hc7,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00B8h] */
                {8'h61,8'hd7,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00BAh] */
                {8'h61,8'hd7,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00BAh] */
                {8'h61,8'he7,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00BCh] */
                {8'h61,8'he7,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00BCh] */
                {8'h61,8'hf7,2'bx0} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00BEh] */
                {8'h61,8'hf7,2'bx1} : dec_cpuwr_enable = 1'b1;  /* CALLT,,[00BEh] */
                {8'h61,8'hcc,2'bx0} : dec_cpuwr_enable = 1'b1;  /* BRK,, */
                {8'h61,8'hcc,2'bx1} : dec_cpuwr_enable = 1'b1;  /* BRK,, */
                {8'h61,8'hdd,2'bxx} : dec_cpuwr_enable = 1'b1;  /* PUSH,,PSW */
                {8'hc1,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* PUSH,,AX */
                {8'hc3,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* PUSH,,BC */
                {8'hc5,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* PUSH,,DE */
                {8'hc7,8'hxx,2'bxx} : dec_cpuwr_enable = 1'b1;  /* PUSH,,HL */
                {8'h31,8'h00,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,saddr.0,$addr8 */
                {8'h31,8'h10,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,saddr.1,$addr8 */
                {8'h31,8'h20,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,saddr.2,$addr8 */
                {8'h31,8'h30,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,saddr.3,$addr8 */
                {8'h31,8'h40,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,saddr.4,$addr8 */
                {8'h31,8'h50,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,saddr.5,$addr8 */
                {8'h31,8'h60,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,saddr.6,$addr8 */
                {8'h31,8'h70,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,saddr.7,$addr8 */
                {8'h31,8'h80,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,sfr.0,$addr8 */
                {8'h31,8'h90,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,sfr.1,$addr8 */
                {8'h31,8'ha0,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,sfr.2,$addr8 */
                {8'h31,8'hb0,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,sfr.3,$addr8 */
                {8'h31,8'hc0,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,sfr.4,$addr8 */
                {8'h31,8'hd0,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,sfr.5,$addr8 */
                {8'h31,8'he0,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,sfr.6,$addr8 */
                {8'h31,8'hf0,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,sfr.7,$addr8 */
                {8'h31,8'h81,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,[HL].0,$addr8 */
                {8'h31,8'h91,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,[HL].1,$addr8 */
                {8'h31,8'ha1,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,[HL].2,$addr8 */
                {8'h31,8'hb1,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,[HL].3,$addr8 */
                {8'h31,8'hc1,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,[HL].4,$addr8 */
                {8'h31,8'hd1,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,[HL].5,$addr8 */
                {8'h31,8'he1,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,[HL].6,$addr8 */
                {8'h31,8'hf1,2'b10} : dec_cpuwr_enable = 1'b1;  /* BTCLR,[HL].7,$addr8 */
                {8'hff,8'hxx,2'bx0} : dec_cpuwr_enable = 1'b1;  /* SOFT,,BREAK */
                {8'hff,8'hxx,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SOFT,,BREAK */
                {8'h61,8'ha1,2'bx0} : dec_cpuwr_enable = 1'b1;  /* SOFT2,,BREAK */
                {8'h61,8'ha1,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SOFT2,,BREAK */
                {8'h61,8'hb1,2'bx0} : dec_cpuwr_enable = 1'b1;  /* SOFT3,,BREAK */
                {8'h61,8'hb1,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SOFT3,,BREAK */
                {8'h61,8'hc1,2'bx0} : dec_cpuwr_enable = 1'b1;  /* SOFT4,,BREAK */
                {8'h61,8'hc1,2'bx1} : dec_cpuwr_enable = 1'b1;  /* SOFT4,,BREAK */
                {8'h61,8'hbb,2'bx1} : dec_cpuwr_enable = 1'b1;  /* XCH,A,sfr */
                {8'h61,8'hba,2'bx1} : dec_cpuwr_enable = 1'b1;  /* XCH,A,!addr16 */
                {8'h61,8'hbe,2'bx1} : dec_cpuwr_enable = 1'b1;  /* XCH,A,[DE] */
                {8'h61,8'hbf,2'bx1} : dec_cpuwr_enable = 1'b1;  /* XCH,A,[DE+byte] */
                {8'h61,8'hbc,2'bx1} : dec_cpuwr_enable = 1'b1;  /* XCH,A,[HL] */
                {8'h61,8'hbd,2'bx1} : dec_cpuwr_enable = 1'b1;  /* XCH,A,[HL+byte] */
                default : dec_cpuwr_enable = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_cpurd_enable;
    reg    dec_cpurd_enable;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 ) begin
            dec_cpurd_enable = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h8d,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV,A,saddr */
                {8'h8e,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV,A,sfr */
                {8'h8f,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV,A,!addr16 */
                {8'h89,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV,A,[DE] */
                {8'h8a,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV,A,[DE+byte] */
                {8'h8b,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV,A,[HL] */
                {8'h8c,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV,A,[HL+byte] */
                {8'h61,8'hc9,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV,A,[HL+B] */
                {8'h61,8'he9,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV,A,[HL+C] */
                {8'h09,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV,A,word[B] */
                {8'h29,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV,A,word[C] */
                {8'h49,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV,A,word[BC] */
                {8'h88,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV,A,[SP+byte] */
                {8'he8,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV,B,saddr */
                {8'he9,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV,B,!addr16 */
                {8'hf8,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV,C,saddr */
                {8'hf9,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV,C,!addr16 */
                {8'hd8,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV,X,saddr */
                {8'hd9,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV,X,!addr16 */
                {8'h61,8'hb8,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV,ES,saddr */
                {8'h61,8'ha8,2'bx0} : dec_cpurd_enable = 1'b1;  /* XCH,A,saddr */
                {8'h61,8'hab,2'bx0} : dec_cpurd_enable = 1'b1;  /* XCH,A,sfr */
                {8'h61,8'haa,2'bx0} : dec_cpurd_enable = 1'b1;  /* XCH,A,!addr16 */
                {8'h61,8'hae,2'bx0} : dec_cpurd_enable = 1'b1;  /* XCH,A,[DE] */
                {8'h61,8'haf,2'bx0} : dec_cpurd_enable = 1'b1;  /* XCH,A,[DE+byte] */
                {8'h61,8'hac,2'bx0} : dec_cpurd_enable = 1'b1;  /* XCH,A,[HL] */
                {8'h61,8'had,2'bx0} : dec_cpurd_enable = 1'b1;  /* XCH,A,[HL+byte] */
                {8'h61,8'hb9,2'bx0} : dec_cpurd_enable = 1'b1;  /* XCH,A,[HL+B] */
                {8'h61,8'ha9,2'bx0} : dec_cpurd_enable = 1'b1;  /* XCH,A,[HL+C] */
                {8'had,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOVW,AX,saddrp */
                {8'hae,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOVW,AX,sfrp */
                {8'haf,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOVW,AX,!addr16 */
                {8'ha9,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOVW,AX,[DE] */
                {8'haa,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOVW,AX,[DE+byte] */
                {8'hab,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOVW,AX,[HL] */
                {8'hac,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOVW,AX,[HL+byte] */
                {8'h59,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOVW,AX,word[B] */
                {8'h69,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOVW,AX,word[C] */
                {8'h79,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOVW,AX,word[BC] */
                {8'ha8,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOVW,AX,[SP+byte] */
                {8'hda,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOVW,BC,saddrp */
                {8'hdb,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOVW,BC,!addr16 */
                {8'hea,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOVW,DE,saddrp */
                {8'heb,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOVW,DE,!addr16 */
                {8'hfa,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOVW,HL,saddrp */
                {8'hfb,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOVW,HL,!addr16 */
                {8'h0a,8'hxx,2'bx0} : dec_cpurd_enable = 1'b1;  /* ADD,saddr,#byte */
                {8'h0b,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* ADD,A,saddr */
                {8'h0f,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* ADD,A,!addr16 */
                {8'h0d,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* ADD,A,[HL] */
                {8'h0e,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* ADD,A,[HL+byte] */
                {8'h61,8'h80,2'bxx} : dec_cpurd_enable = 1'b1;  /* ADD,A,[HL+B] */
                {8'h61,8'h82,2'bxx} : dec_cpurd_enable = 1'b1;  /* ADD,A,[HL+C] */
                {8'h1a,8'hxx,2'bx0} : dec_cpurd_enable = 1'b1;  /* ADDC,saddr,#byte */
                {8'h1b,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* ADDC,A,saddr */
                {8'h1f,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* ADDC,A,!addr16 */
                {8'h1d,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* ADDC,A,[HL] */
                {8'h1e,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* ADDC,A,[HL+byte] */
                {8'h61,8'h90,2'bxx} : dec_cpurd_enable = 1'b1;  /* ADDC,A,[HL+B] */
                {8'h61,8'h92,2'bxx} : dec_cpurd_enable = 1'b1;  /* ADDC,A,[HL+C] */
                {8'h2a,8'hxx,2'bx0} : dec_cpurd_enable = 1'b1;  /* SUB,saddr,#byte */
                {8'h2b,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* SUB,A,saddr */
                {8'h2f,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* SUB,A,!addr16 */
                {8'h2d,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* SUB,A,[HL] */
                {8'h2e,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* SUB,A,[HL+byte] */
                {8'h61,8'ha0,2'bxx} : dec_cpurd_enable = 1'b1;  /* SUB,A,[HL+B] */
                {8'h61,8'ha2,2'bxx} : dec_cpurd_enable = 1'b1;  /* SUB,A,[HL+C] */
                {8'h3a,8'hxx,2'bx0} : dec_cpurd_enable = 1'b1;  /* SUBC,saddr,#byte */
                {8'h3b,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* SUBC,A,saddr */
                {8'h3f,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* SUBC,A,!addr16 */
                {8'h3d,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* SUBC,A,[HL] */
                {8'h3e,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* SUBC,A,[HL+byte] */
                {8'h61,8'hb0,2'bxx} : dec_cpurd_enable = 1'b1;  /* SUBC,A,[HL+B] */
                {8'h61,8'hb2,2'bxx} : dec_cpurd_enable = 1'b1;  /* SUBC,A,[HL+C] */
                {8'h5a,8'hxx,2'bx0} : dec_cpurd_enable = 1'b1;  /* AND,saddr,#byte */
                {8'h5b,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND,A,saddr */
                {8'h5f,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND,A,!addr16 */
                {8'h5d,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND,A,[HL] */
                {8'h5e,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND,A,[HL+byte] */
                {8'h61,8'hd0,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND,A,[HL+B] */
                {8'h61,8'hd2,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND,A,[HL+C] */
                {8'h6a,8'hxx,2'bx0} : dec_cpurd_enable = 1'b1;  /* OR,saddr,#byte */
                {8'h6b,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR,A,saddr */
                {8'h6f,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR,A,!addr16 */
                {8'h6d,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR,A,[HL] */
                {8'h6e,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR,A,[HL+byte] */
                {8'h61,8'he0,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR,A,[HL+B] */
                {8'h61,8'he2,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR,A,[HL+C] */
                {8'h7a,8'hxx,2'bx0} : dec_cpurd_enable = 1'b1;  /* XOR,saddr,#byte */
                {8'h7b,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR,A,saddr */
                {8'h7f,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR,A,!addr16 */
                {8'h7d,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR,A,[HL] */
                {8'h7e,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR,A,[HL+byte] */
                {8'h61,8'hf0,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR,A,[HL+B] */
                {8'h61,8'hf2,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR,A,[HL+C] */
                {8'h4a,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* CMP,saddr,#byte */
                {8'h40,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* CMP,!addr16,#byte */
                {8'h4b,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* CMP,A,saddr */
                {8'h4f,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* CMP,A,!addr16 */
                {8'h4d,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* CMP,A,[HL] */
                {8'h4e,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* CMP,A,[HL+byte] */
                {8'h61,8'hc0,2'bxx} : dec_cpurd_enable = 1'b1;  /* CMP,A,[HL+B] */
                {8'h61,8'hc2,2'bxx} : dec_cpurd_enable = 1'b1;  /* CMP,A,[HL+C] */
                {8'h61,8'hde,2'bxx} : dec_cpurd_enable = 1'b1;  /* CMPS,X,[HL+byte] */
                {8'hd4,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* CMP0,,saddr */
                {8'hd5,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* CMP0,,!addr16 */
                {8'h06,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* ADDW,AX,saddrp */
                {8'h02,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* ADDW,AX,!addr16 */
                {8'h61,8'h09,2'bxx} : dec_cpurd_enable = 1'b1;  /* ADDW,AX,[HL+byte] */
                {8'h26,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* SUBW,AX,saddrp */
                {8'h22,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* SUBW,AX,!addr16 */
                {8'h61,8'h29,2'bxx} : dec_cpurd_enable = 1'b1;  /* SUBW,AX,[HL+byte] */
                {8'h46,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* CMPW,AX,saddrp */
                {8'h42,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* CMPW,AX,!addr16 */
                {8'h61,8'h49,2'bxx} : dec_cpurd_enable = 1'b1;  /* CMPW,AX,[HL+byte] */
                {8'ha4,8'hxx,2'bx0} : dec_cpurd_enable = 1'b1;  /* INC,,saddr */
                {8'ha0,8'hxx,2'bx0} : dec_cpurd_enable = 1'b1;  /* INC,,!addr16 */
                {8'h61,8'h59,2'bx0} : dec_cpurd_enable = 1'b1;  /* INC,,[HL+byte] */
                {8'hb4,8'hxx,2'bx0} : dec_cpurd_enable = 1'b1;  /* DEC,,saddr */
                {8'hb0,8'hxx,2'bx0} : dec_cpurd_enable = 1'b1;  /* DEC,,!addr16 */
                {8'h61,8'h69,2'bx0} : dec_cpurd_enable = 1'b1;  /* DEC,,[HL+byte] */
                {8'ha6,8'hxx,2'bx0} : dec_cpurd_enable = 1'b1;  /* INCW,,saddrp */
                {8'ha2,8'hxx,2'bx0} : dec_cpurd_enable = 1'b1;  /* INCW,,!addr16 */
                {8'h61,8'h79,2'bx0} : dec_cpurd_enable = 1'b1;  /* INCW,,[HL+byte] */
                {8'hb6,8'hxx,2'bx0} : dec_cpurd_enable = 1'b1;  /* DECW,,saddrp */
                {8'hb2,8'hxx,2'bx0} : dec_cpurd_enable = 1'b1;  /* DECW,,!addr16 */
                {8'h61,8'h89,2'bx0} : dec_cpurd_enable = 1'b1;  /* DECW,,[HL+byte] */
                {8'h71,8'h04,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,saddr.0 */
                {8'h71,8'h14,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,saddr.1 */
                {8'h71,8'h24,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,saddr.2 */
                {8'h71,8'h34,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,saddr.3 */
                {8'h71,8'h44,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,saddr.4 */
                {8'h71,8'h54,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,saddr.5 */
                {8'h71,8'h64,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,saddr.6 */
                {8'h71,8'h74,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,saddr.7 */
                {8'h71,8'h0c,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,sfr.0 */
                {8'h71,8'h1c,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,sfr.1 */
                {8'h71,8'h2c,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,sfr.2 */
                {8'h71,8'h3c,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,sfr.3 */
                {8'h71,8'h4c,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,sfr.4 */
                {8'h71,8'h5c,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,sfr.5 */
                {8'h71,8'h6c,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,sfr.6 */
                {8'h71,8'h7c,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,sfr.7 */
                {8'h71,8'h84,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,[HL].0 */
                {8'h71,8'h94,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,[HL].1 */
                {8'h71,8'ha4,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,[HL].2 */
                {8'h71,8'hb4,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,[HL].3 */
                {8'h71,8'hc4,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,[HL].4 */
                {8'h71,8'hd4,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,[HL].5 */
                {8'h71,8'he4,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,[HL].6 */
                {8'h71,8'hf4,2'bxx} : dec_cpurd_enable = 1'b1;  /* MOV1,CY,[HL].7 */
                {8'h71,8'h01,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,saddr.0,CY */
                {8'h71,8'h11,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,saddr.1,CY */
                {8'h71,8'h21,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,saddr.2,CY */
                {8'h71,8'h31,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,saddr.3,CY */
                {8'h71,8'h41,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,saddr.4,CY */
                {8'h71,8'h51,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,saddr.5,CY */
                {8'h71,8'h61,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,saddr.6,CY */
                {8'h71,8'h71,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,saddr.7,CY */
                {8'h71,8'h09,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,sfr.0,CY */
                {8'h71,8'h19,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,sfr.1,CY */
                {8'h71,8'h29,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,sfr.2,CY */
                {8'h71,8'h39,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,sfr.3,CY */
                {8'h71,8'h49,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,sfr.4,CY */
                {8'h71,8'h59,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,sfr.5,CY */
                {8'h71,8'h69,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,sfr.6,CY */
                {8'h71,8'h79,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,sfr.7,CY */
                {8'h71,8'h81,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,[HL].0,CY */
                {8'h71,8'h91,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,[HL].1,CY */
                {8'h71,8'ha1,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,[HL].2,CY */
                {8'h71,8'hb1,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,[HL].3,CY */
                {8'h71,8'hc1,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,[HL].4,CY */
                {8'h71,8'hd1,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,[HL].5,CY */
                {8'h71,8'he1,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,[HL].6,CY */
                {8'h71,8'hf1,2'bx0} : dec_cpurd_enable = 1'b1;  /* MOV1,[HL].7,CY */
                {8'h71,8'h05,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,saddr.0 */
                {8'h71,8'h15,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,saddr.1 */
                {8'h71,8'h25,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,saddr.2 */
                {8'h71,8'h35,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,saddr.3 */
                {8'h71,8'h45,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,saddr.4 */
                {8'h71,8'h55,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,saddr.5 */
                {8'h71,8'h65,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,saddr.6 */
                {8'h71,8'h75,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,saddr.7 */
                {8'h71,8'h0d,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,sfr.0 */
                {8'h71,8'h1d,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,sfr.1 */
                {8'h71,8'h2d,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,sfr.2 */
                {8'h71,8'h3d,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,sfr.3 */
                {8'h71,8'h4d,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,sfr.4 */
                {8'h71,8'h5d,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,sfr.5 */
                {8'h71,8'h6d,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,sfr.6 */
                {8'h71,8'h7d,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,sfr.7 */
                {8'h71,8'h85,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,[HL].0 */
                {8'h71,8'h95,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,[HL].1 */
                {8'h71,8'ha5,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,[HL].2 */
                {8'h71,8'hb5,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,[HL].3 */
                {8'h71,8'hc5,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,[HL].4 */
                {8'h71,8'hd5,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,[HL].5 */
                {8'h71,8'he5,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,[HL].6 */
                {8'h71,8'hf5,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND1,CY,[HL].7 */
                {8'h71,8'h06,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,saddr.0 */
                {8'h71,8'h16,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,saddr.1 */
                {8'h71,8'h26,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,saddr.2 */
                {8'h71,8'h36,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,saddr.3 */
                {8'h71,8'h46,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,saddr.4 */
                {8'h71,8'h56,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,saddr.5 */
                {8'h71,8'h66,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,saddr.6 */
                {8'h71,8'h76,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,saddr.7 */
                {8'h71,8'h0e,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,sfr.0 */
                {8'h71,8'h1e,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,sfr.1 */
                {8'h71,8'h2e,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,sfr.2 */
                {8'h71,8'h3e,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,sfr.3 */
                {8'h71,8'h4e,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,sfr.4 */
                {8'h71,8'h5e,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,sfr.5 */
                {8'h71,8'h6e,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,sfr.6 */
                {8'h71,8'h7e,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,sfr.7 */
                {8'h71,8'h86,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,[HL].0 */
                {8'h71,8'h96,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,[HL].1 */
                {8'h71,8'ha6,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,[HL].2 */
                {8'h71,8'hb6,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,[HL].3 */
                {8'h71,8'hc6,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,[HL].4 */
                {8'h71,8'hd6,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,[HL].5 */
                {8'h71,8'he6,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,[HL].6 */
                {8'h71,8'hf6,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR1,CY,[HL].7 */
                {8'h71,8'h07,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,saddr.0 */
                {8'h71,8'h17,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,saddr.1 */
                {8'h71,8'h27,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,saddr.2 */
                {8'h71,8'h37,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,saddr.3 */
                {8'h71,8'h47,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,saddr.4 */
                {8'h71,8'h57,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,saddr.5 */
                {8'h71,8'h67,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,saddr.6 */
                {8'h71,8'h77,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,saddr.7 */
                {8'h71,8'h0f,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,sfr.0 */
                {8'h71,8'h1f,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,sfr.1 */
                {8'h71,8'h2f,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,sfr.2 */
                {8'h71,8'h3f,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,sfr.3 */
                {8'h71,8'h4f,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,sfr.4 */
                {8'h71,8'h5f,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,sfr.5 */
                {8'h71,8'h6f,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,sfr.6 */
                {8'h71,8'h7f,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,sfr.7 */
                {8'h71,8'h87,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,[HL].0 */
                {8'h71,8'h97,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,[HL].1 */
                {8'h71,8'ha7,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,[HL].2 */
                {8'h71,8'hb7,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,[HL].3 */
                {8'h71,8'hc7,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,[HL].4 */
                {8'h71,8'hd7,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,[HL].5 */
                {8'h71,8'he7,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,[HL].6 */
                {8'h71,8'hf7,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR1,CY,[HL].7 */
                {8'h71,8'h02,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,saddr.0 */
                {8'h71,8'h12,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,saddr.1 */
                {8'h71,8'h22,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,saddr.2 */
                {8'h71,8'h32,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,saddr.3 */
                {8'h71,8'h42,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,saddr.4 */
                {8'h71,8'h52,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,saddr.5 */
                {8'h71,8'h62,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,saddr.6 */
                {8'h71,8'h72,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,saddr.7 */
                {8'h71,8'h0a,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,sfr.0 */
                {8'h71,8'h1a,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,sfr.1 */
                {8'h71,8'h2a,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,sfr.2 */
                {8'h71,8'h3a,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,sfr.3 */
                {8'h71,8'h4a,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,sfr.4 */
                {8'h71,8'h5a,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,sfr.5 */
                {8'h71,8'h6a,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,sfr.6 */
                {8'h71,8'h7a,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,sfr.7 */
                {8'h71,8'h00,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,!addr16.0 */
                {8'h71,8'h10,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,!addr16.1 */
                {8'h71,8'h20,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,!addr16.2 */
                {8'h71,8'h30,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,!addr16.3 */
                {8'h71,8'h40,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,!addr16.4 */
                {8'h71,8'h50,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,!addr16.5 */
                {8'h71,8'h60,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,!addr16.6 */
                {8'h71,8'h70,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,!addr16.7 */
                {8'h71,8'h82,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,[HL].0 */
                {8'h71,8'h92,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,[HL].1 */
                {8'h71,8'ha2,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,[HL].2 */
                {8'h71,8'hb2,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,[HL].3 */
                {8'h71,8'hc2,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,[HL].4 */
                {8'h71,8'hd2,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,[HL].5 */
                {8'h71,8'he2,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,[HL].6 */
                {8'h71,8'hf2,2'bx0} : dec_cpurd_enable = 1'b1;  /* SET1,,[HL].7 */
                {8'h71,8'h03,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,saddr.0 */
                {8'h71,8'h13,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,saddr.1 */
                {8'h71,8'h23,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,saddr.2 */
                {8'h71,8'h33,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,saddr.3 */
                {8'h71,8'h43,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,saddr.4 */
                {8'h71,8'h53,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,saddr.5 */
                {8'h71,8'h63,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,saddr.6 */
                {8'h71,8'h73,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,saddr.7 */
                {8'h71,8'h0b,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,sfr.0 */
                {8'h71,8'h1b,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,sfr.1 */
                {8'h71,8'h2b,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,sfr.2 */
                {8'h71,8'h3b,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,sfr.3 */
                {8'h71,8'h4b,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,sfr.4 */
                {8'h71,8'h5b,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,sfr.5 */
                {8'h71,8'h6b,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,sfr.6 */
                {8'h71,8'h7b,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,sfr.7 */
                {8'h71,8'h08,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,!addr16.0 */
                {8'h71,8'h18,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,!addr16.1 */
                {8'h71,8'h28,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,!addr16.2 */
                {8'h71,8'h38,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,!addr16.3 */
                {8'h71,8'h48,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,!addr16.4 */
                {8'h71,8'h58,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,!addr16.5 */
                {8'h71,8'h68,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,!addr16.6 */
                {8'h71,8'h78,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,!addr16.7 */
                {8'h71,8'h83,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,[HL].0 */
                {8'h71,8'h93,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,[HL].1 */
                {8'h71,8'ha3,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,[HL].2 */
                {8'h71,8'hb3,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,[HL].3 */
                {8'h71,8'hc3,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,[HL].4 */
                {8'h71,8'hd3,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,[HL].5 */
                {8'h71,8'he3,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,[HL].6 */
                {8'h71,8'hf3,2'bx0} : dec_cpurd_enable = 1'b1;  /* CLR1,,[HL].7 */
                {8'hd7,8'hxx,2'b00} : dec_cpurd_enable = 1'b1;  /* RET,, */
                {8'hd7,8'hxx,2'b01} : dec_cpurd_enable = 1'b1;  /* RET,, */
                {8'h61,8'hec,2'b00} : dec_cpurd_enable = 1'b1;  /* RETB,, */
                {8'h61,8'hec,2'b01} : dec_cpurd_enable = 1'b1;  /* RETB,, */
                {8'h61,8'hfc,2'b00} : dec_cpurd_enable = 1'b1;  /* RETI,, */
                {8'h61,8'hfc,2'b01} : dec_cpurd_enable = 1'b1;  /* RETI,, */
                {8'h61,8'hcd,2'bxx} : dec_cpurd_enable = 1'b1;  /* POP,,PSW */
                {8'hc0,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* POP,,AX */
                {8'hc2,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* POP,,BC */
                {8'hc4,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* POP,,DE */
                {8'hc6,8'hxx,2'bxx} : dec_cpurd_enable = 1'b1;  /* POP,,HL */
                {8'h31,8'h02,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,saddr.0,$addr8 */
                {8'h31,8'h12,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,saddr.1,$addr8 */
                {8'h31,8'h22,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,saddr.2,$addr8 */
                {8'h31,8'h32,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,saddr.3,$addr8 */
                {8'h31,8'h42,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,saddr.4,$addr8 */
                {8'h31,8'h52,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,saddr.5,$addr8 */
                {8'h31,8'h62,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,saddr.6,$addr8 */
                {8'h31,8'h72,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,saddr.7,$addr8 */
                {8'h31,8'h82,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,sfr.0,$addr8 */
                {8'h31,8'h92,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,sfr.1,$addr8 */
                {8'h31,8'ha2,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,sfr.2,$addr8 */
                {8'h31,8'hb2,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,sfr.3,$addr8 */
                {8'h31,8'hc2,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,sfr.4,$addr8 */
                {8'h31,8'hd2,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,sfr.5,$addr8 */
                {8'h31,8'he2,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,sfr.6,$addr8 */
                {8'h31,8'hf2,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,sfr.7,$addr8 */
                {8'h31,8'h83,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,[HL].0,$addr8 */
                {8'h31,8'h93,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,[HL].1,$addr8 */
                {8'h31,8'ha3,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,[HL].2,$addr8 */
                {8'h31,8'hb3,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,[HL].3,$addr8 */
                {8'h31,8'hc3,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,[HL].4,$addr8 */
                {8'h31,8'hd3,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,[HL].5,$addr8 */
                {8'h31,8'he3,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,[HL].6,$addr8 */
                {8'h31,8'hf3,2'b00} : dec_cpurd_enable = 1'b1;  /* BT,[HL].7,$addr8 */
                {8'h31,8'h04,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,saddr.0,$addr8 */
                {8'h31,8'h14,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,saddr.1,$addr8 */
                {8'h31,8'h24,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,saddr.2,$addr8 */
                {8'h31,8'h34,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,saddr.3,$addr8 */
                {8'h31,8'h44,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,saddr.4,$addr8 */
                {8'h31,8'h54,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,saddr.5,$addr8 */
                {8'h31,8'h64,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,saddr.6,$addr8 */
                {8'h31,8'h74,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,saddr.7,$addr8 */
                {8'h31,8'h84,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,sfr.0,$addr8 */
                {8'h31,8'h94,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,sfr.1,$addr8 */
                {8'h31,8'ha4,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,sfr.2,$addr8 */
                {8'h31,8'hb4,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,sfr.3,$addr8 */
                {8'h31,8'hc4,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,sfr.4,$addr8 */
                {8'h31,8'hd4,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,sfr.5,$addr8 */
                {8'h31,8'he4,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,sfr.6,$addr8 */
                {8'h31,8'hf4,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,sfr.7,$addr8 */
                {8'h31,8'h85,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,[HL].0,$addr8 */
                {8'h31,8'h95,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,[HL].1,$addr8 */
                {8'h31,8'ha5,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,[HL].2,$addr8 */
                {8'h31,8'hb5,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,[HL].3,$addr8 */
                {8'h31,8'hc5,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,[HL].4,$addr8 */
                {8'h31,8'hd5,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,[HL].5,$addr8 */
                {8'h31,8'he5,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,[HL].6,$addr8 */
                {8'h31,8'hf5,2'b00} : dec_cpurd_enable = 1'b1;  /* BF,[HL].7,$addr8 */
                {8'h31,8'h00,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,saddr.0,$addr8 */
                {8'h31,8'h00,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,saddr.0,$addr8 */
                {8'h31,8'h10,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,saddr.1,$addr8 */
                {8'h31,8'h10,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,saddr.1,$addr8 */
                {8'h31,8'h20,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,saddr.2,$addr8 */
                {8'h31,8'h20,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,saddr.2,$addr8 */
                {8'h31,8'h30,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,saddr.3,$addr8 */
                {8'h31,8'h30,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,saddr.3,$addr8 */
                {8'h31,8'h40,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,saddr.4,$addr8 */
                {8'h31,8'h40,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,saddr.4,$addr8 */
                {8'h31,8'h50,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,saddr.5,$addr8 */
                {8'h31,8'h50,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,saddr.5,$addr8 */
                {8'h31,8'h60,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,saddr.6,$addr8 */
                {8'h31,8'h60,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,saddr.6,$addr8 */
                {8'h31,8'h70,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,saddr.7,$addr8 */
                {8'h31,8'h70,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,saddr.7,$addr8 */
                {8'h31,8'h80,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,sfr.0,$addr8 */
                {8'h31,8'h80,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,sfr.0,$addr8 */
                {8'h31,8'h90,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,sfr.1,$addr8 */
                {8'h31,8'h90,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,sfr.1,$addr8 */
                {8'h31,8'ha0,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,sfr.2,$addr8 */
                {8'h31,8'ha0,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,sfr.2,$addr8 */
                {8'h31,8'hb0,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,sfr.3,$addr8 */
                {8'h31,8'hb0,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,sfr.3,$addr8 */
                {8'h31,8'hc0,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,sfr.4,$addr8 */
                {8'h31,8'hc0,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,sfr.4,$addr8 */
                {8'h31,8'hd0,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,sfr.5,$addr8 */
                {8'h31,8'hd0,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,sfr.5,$addr8 */
                {8'h31,8'he0,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,sfr.6,$addr8 */
                {8'h31,8'he0,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,sfr.6,$addr8 */
                {8'h31,8'hf0,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,sfr.7,$addr8 */
                {8'h31,8'hf0,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,sfr.7,$addr8 */
                {8'h31,8'h81,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,[HL].0,$addr8 */
                {8'h31,8'h81,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,[HL].0,$addr8 */
                {8'h31,8'h91,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,[HL].1,$addr8 */
                {8'h31,8'h91,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,[HL].1,$addr8 */
                {8'h31,8'ha1,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,[HL].2,$addr8 */
                {8'h31,8'ha1,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,[HL].2,$addr8 */
                {8'h31,8'hb1,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,[HL].3,$addr8 */
                {8'h31,8'hb1,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,[HL].3,$addr8 */
                {8'h31,8'hc1,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,[HL].4,$addr8 */
                {8'h31,8'hc1,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,[HL].4,$addr8 */
                {8'h31,8'hd1,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,[HL].5,$addr8 */
                {8'h31,8'hd1,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,[HL].5,$addr8 */
                {8'h31,8'he1,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,[HL].6,$addr8 */
                {8'h31,8'he1,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,[HL].6,$addr8 */
                {8'h31,8'hf1,2'b00} : dec_cpurd_enable = 1'b1;  /* BTCLR,[HL].7,$addr8 */
                {8'h31,8'hf1,2'b01} : dec_cpurd_enable = 1'b1;  /* BTCLR,[HL].7,$addr8 */
                {8'h61,8'hbb,2'bx0} : dec_cpurd_enable = 1'b1;  /* XCH,A,sfr */
                {8'h61,8'hba,2'bx0} : dec_cpurd_enable = 1'b1;  /* XCH,A,!addr16 */
                {8'h61,8'hbe,2'bx0} : dec_cpurd_enable = 1'b1;  /* XCH,A,[DE] */
                {8'h61,8'hbf,2'bx0} : dec_cpurd_enable = 1'b1;  /* XCH,A,[DE+byte] */
                {8'h61,8'hbc,2'bx0} : dec_cpurd_enable = 1'b1;  /* XCH,A,[HL] */
                {8'h61,8'hbd,2'bx0} : dec_cpurd_enable = 1'b1;  /* XCH,A,[HL+byte] */
                {8'h61,8'hd1,2'bxx} : dec_cpurd_enable = 1'b1;  /* AND,A,[HL+B] */
                {8'h61,8'he1,2'bxx} : dec_cpurd_enable = 1'b1;  /* OR,A,[HL+B] */
                {8'h61,8'hf1,2'bxx} : dec_cpurd_enable = 1'b1;  /* XOR,A,[HL+B] */
                {8'h61,8'h83,2'bxx} : dec_cpurd_enable = 1'b1;  /* ADD,A,[HL+C] */
                {8'h61,8'h93,2'bxx} : dec_cpurd_enable = 1'b1;  /* ADDC,A,[HL+C] */
                {8'h61,8'ha3,2'bxx} : dec_cpurd_enable = 1'b1;  /* SUB,A,[HL+C] */
                {8'h61,8'hb3,2'bxx} : dec_cpurd_enable = 1'b1;  /* SUBC,A,[HL+C] */
                default : dec_cpurd_enable = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ma_enable;
    reg    dec_ma_enable;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(decout_mask == 1'b1) begin
//            dec_ma_enable = 1'b0;
//        end else if(rstvec == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1) begin
            dec_ma_enable = 1'b0;
        end else if(ivack == 1'b1) begin
            casex ({stage_adr})  
                {2'b00} : dec_ma_enable = 1'b1;  /* Interrupt */
                {2'b01} : dec_ma_enable = 1'b1;  /* Interrupt */
                default : dec_ma_enable = 1'b0;
            endcase
        end else if(skpack == 1'b1) begin
            dec_ma_enable = 1'b0;
        end else begin
            if(ID_stage0 == 8'h61) begin
                casex ({ID_stage1,stage_adr})  
                    {8'hc9,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,A,[HL+B] */
                    {8'hd9,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,[HL+B],A */
                    {8'he9,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,A,[HL+C] */
                    {8'hf9,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,[HL+C],A */
                    {8'hb8,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,ES,saddr */
                    {8'hce,2'bxx} : dec_ma_enable = 1'b1;  /* MOVS,[HL+byte],X */
                    {8'ha8,2'bx0} : dec_ma_enable = 1'b1;  /* XCH,A,saddr */
                    {8'ha8,2'bx1} : dec_ma_enable = 1'b1;  /* XCH,A,saddr */
                    {8'hab,2'bx0} : dec_ma_enable = 1'b1;  /* XCH,A,sfr */
                    {8'hab,2'bx1} : dec_ma_enable = 1'b1;  /* XCH,A,sfr */
                    {8'haa,2'bx0} : dec_ma_enable = 1'b1;  /* XCH,A,!addr16 */
                    {8'haa,2'bx1} : dec_ma_enable = 1'b1;  /* XCH,A,!addr16 */
                    {8'hae,2'bx0} : dec_ma_enable = 1'b1;  /* XCH,A,[DE] */
                    {8'hae,2'bx1} : dec_ma_enable = 1'b1;  /* XCH,A,[DE] */
                    {8'haf,2'bx0} : dec_ma_enable = 1'b1;  /* XCH,A,[DE+byte] */
                    {8'haf,2'bx1} : dec_ma_enable = 1'b1;  /* XCH,A,[DE+byte] */
                    {8'hac,2'bx0} : dec_ma_enable = 1'b1;  /* XCH,A,[HL] */
                    {8'hac,2'bx1} : dec_ma_enable = 1'b1;  /* XCH,A,[HL] */
                    {8'had,2'bx0} : dec_ma_enable = 1'b1;  /* XCH,A,[HL+byte] */
                    {8'had,2'bx1} : dec_ma_enable = 1'b1;  /* XCH,A,[HL+byte] */
                    {8'hb9,2'bx0} : dec_ma_enable = 1'b1;  /* XCH,A,[HL+B] */
                    {8'hb9,2'bx1} : dec_ma_enable = 1'b1;  /* XCH,A,[HL+B] */
                    {8'ha9,2'bx0} : dec_ma_enable = 1'b1;  /* XCH,A,[HL+C] */
                    {8'ha9,2'bx1} : dec_ma_enable = 1'b1;  /* XCH,A,[HL+C] */
                    {8'h80,2'bxx} : dec_ma_enable = 1'b1;  /* ADD,A,[HL+B] */
                    {8'h82,2'bxx} : dec_ma_enable = 1'b1;  /* ADD,A,[HL+C] */
                    {8'h90,2'bxx} : dec_ma_enable = 1'b1;  /* ADDC,A,[HL+B] */
                    {8'h92,2'bxx} : dec_ma_enable = 1'b1;  /* ADDC,A,[HL+C] */
                    {8'ha0,2'bxx} : dec_ma_enable = 1'b1;  /* SUB,A,[HL+B] */
                    {8'ha2,2'bxx} : dec_ma_enable = 1'b1;  /* SUB,A,[HL+C] */
                    {8'hb0,2'bxx} : dec_ma_enable = 1'b1;  /* SUBC,A,[HL+B] */
                    {8'hb2,2'bxx} : dec_ma_enable = 1'b1;  /* SUBC,A,[HL+C] */
                    {8'hd0,2'bxx} : dec_ma_enable = 1'b1;  /* AND,A,[HL+B] */
                    {8'hd2,2'bxx} : dec_ma_enable = 1'b1;  /* AND,A,[HL+C] */
                    {8'he0,2'bxx} : dec_ma_enable = 1'b1;  /* OR,A,[HL+B] */
                    {8'he2,2'bxx} : dec_ma_enable = 1'b1;  /* OR,A,[HL+C] */
                    {8'hf0,2'bxx} : dec_ma_enable = 1'b1;  /* XOR,A,[HL+B] */
                    {8'hf2,2'bxx} : dec_ma_enable = 1'b1;  /* XOR,A,[HL+C] */
                    {8'hc0,2'bxx} : dec_ma_enable = 1'b1;  /* CMP,A,[HL+B] */
                    {8'hc2,2'bxx} : dec_ma_enable = 1'b1;  /* CMP,A,[HL+C] */
                    {8'hde,2'bxx} : dec_ma_enable = 1'b1;  /* CMPS,X,[HL+byte] */
                    {8'h09,2'bxx} : dec_ma_enable = 1'b1;  /* ADDW,AX,[HL+byte] */
                    {8'h29,2'bxx} : dec_ma_enable = 1'b1;  /* SUBW,AX,[HL+byte] */
                    {8'h49,2'bxx} : dec_ma_enable = 1'b1;  /* CMPW,AX,[HL+byte] */
                    {8'h59,2'bx0} : dec_ma_enable = 1'b1;  /* INC,,[HL+byte] */
                    {8'h59,2'bx1} : dec_ma_enable = 1'b1;  /* INC,,[HL+byte] */
                    {8'h69,2'bx0} : dec_ma_enable = 1'b1;  /* DEC,,[HL+byte] */
                    {8'h69,2'bx1} : dec_ma_enable = 1'b1;  /* DEC,,[HL+byte] */
                    {8'h79,2'bx0} : dec_ma_enable = 1'b1;  /* INCW,,[HL+byte] */
                    {8'h79,2'bx1} : dec_ma_enable = 1'b1;  /* INCW,,[HL+byte] */
                    {8'h89,2'bx0} : dec_ma_enable = 1'b1;  /* DECW,,[HL+byte] */
                    {8'h89,2'bx1} : dec_ma_enable = 1'b1;  /* DECW,,[HL+byte] */
                    {8'hca,2'bx0} : dec_ma_enable = 1'b1;  /* CALL,,AX */
                    {8'hca,2'bx1} : dec_ma_enable = 1'b1;  /* CALL,,AX */
                    {8'hda,2'bx0} : dec_ma_enable = 1'b1;  /* CALL,,BC */
                    {8'hda,2'bx1} : dec_ma_enable = 1'b1;  /* CALL,,BC */
                    {8'hea,2'bx0} : dec_ma_enable = 1'b1;  /* CALL,,DE */
                    {8'hea,2'bx1} : dec_ma_enable = 1'b1;  /* CALL,,DE */
                    {8'hfa,2'bx0} : dec_ma_enable = 1'b1;  /* CALL,,HL */
                    {8'hfa,2'bx1} : dec_ma_enable = 1'b1;  /* CALL,,HL */
                    {8'h84,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[0080h] */
                    {8'h84,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[0080h] */
                    {8'h94,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[0082h] */
                    {8'h94,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[0082h] */
                    {8'ha4,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[0084h] */
                    {8'ha4,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[0084h] */
                    {8'hb4,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[0086h] */
                    {8'hb4,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[0086h] */
                    {8'hc4,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[0088h] */
                    {8'hc4,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[0088h] */
                    {8'hd4,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[008Ah] */
                    {8'hd4,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[008Ah] */
                    {8'he4,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[008Ch] */
                    {8'he4,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[008Ch] */
                    {8'hf4,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[008Eh] */
                    {8'hf4,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[008Eh] */
                    {8'h85,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[0090h] */
                    {8'h85,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[0090h] */
                    {8'h95,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[0092h] */
                    {8'h95,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[0092h] */
                    {8'ha5,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[0094h] */
                    {8'ha5,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[0094h] */
                    {8'hb5,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[0096h] */
                    {8'hb5,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[0096h] */
                    {8'hc5,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[0098h] */
                    {8'hc5,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[0098h] */
                    {8'hd5,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[009Ah] */
                    {8'hd5,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[009Ah] */
                    {8'he5,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[009Ch] */
                    {8'he5,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[009Ch] */
                    {8'hf5,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[009Eh] */
                    {8'hf5,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[009Eh] */
                    {8'h86,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[00A0h] */
                    {8'h86,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[00A0h] */
                    {8'h96,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[00A2h] */
                    {8'h96,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[00A2h] */
                    {8'ha6,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[00A4h] */
                    {8'ha6,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[00A4h] */
                    {8'hb6,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[00A6h] */
                    {8'hb6,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[00A6h] */
                    {8'hc6,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[00A8h] */
                    {8'hc6,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[00A8h] */
                    {8'hd6,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[00AAh] */
                    {8'hd6,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[00AAh] */
                    {8'he6,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[00ACh] */
                    {8'he6,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[00ACh] */
                    {8'hf6,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[00AEh] */
                    {8'hf6,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[00AEh] */
                    {8'h87,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[00B0h] */
                    {8'h87,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[00B0h] */
                    {8'h97,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[00B2h] */
                    {8'h97,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[00B2h] */
                    {8'ha7,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[00B4h] */
                    {8'ha7,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[00B4h] */
                    {8'hb7,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[00B6h] */
                    {8'hb7,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[00B6h] */
                    {8'hc7,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[00B8h] */
                    {8'hc7,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[00B8h] */
                    {8'hd7,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[00BAh] */
                    {8'hd7,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[00BAh] */
                    {8'he7,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[00BCh] */
                    {8'he7,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[00BCh] */
                    {8'hf7,2'bx0} : dec_ma_enable = 1'b1;  /* CALLT,,[00BEh] */
                    {8'hf7,2'bx1} : dec_ma_enable = 1'b1;  /* CALLT,,[00BEh] */
                    {8'hcc,2'bx0} : dec_ma_enable = 1'b1;  /* BRK,, */
                    {8'hcc,2'bx1} : dec_ma_enable = 1'b1;  /* BRK,, */
                    {8'hec,2'b00} : dec_ma_enable = 1'b1;  /* RETB,, */
                    {8'hec,2'b01} : dec_ma_enable = 1'b1;  /* RETB,, */
                    {8'hfc,2'b00} : dec_ma_enable = 1'b1;  /* RETI,, */
                    {8'hfc,2'b01} : dec_ma_enable = 1'b1;  /* RETI,, */
                    {8'hdd,2'bxx} : dec_ma_enable = 1'b1;  /* PUSH,,PSW */
                    {8'hcd,2'bxx} : dec_ma_enable = 1'b1;  /* POP,,PSW */
                    {8'ha1,2'bx0} : dec_ma_enable = 1'b1;  /* SOFT2,,BREAK */
                    {8'ha1,2'bx1} : dec_ma_enable = 1'b1;  /* SOFT2,,BREAK */
                    {8'hb1,2'bx0} : dec_ma_enable = 1'b1;  /* SOFT3,,BREAK */
                    {8'hb1,2'bx1} : dec_ma_enable = 1'b1;  /* SOFT3,,BREAK */
                    {8'hc1,2'bx0} : dec_ma_enable = 1'b1;  /* SOFT4,,BREAK */
                    {8'hc1,2'bx1} : dec_ma_enable = 1'b1;  /* SOFT4,,BREAK */
                    {8'hbb,2'bx0} : dec_ma_enable = 1'b1;  /* XCH,A,sfr */
                    {8'hbb,2'bx1} : dec_ma_enable = 1'b1;  /* XCH,A,sfr */
                    {8'hba,2'bx0} : dec_ma_enable = 1'b1;  /* XCH,A,!addr16 */
                    {8'hba,2'bx1} : dec_ma_enable = 1'b1;  /* XCH,A,!addr16 */
                    {8'hbe,2'bx0} : dec_ma_enable = 1'b1;  /* XCH,A,[DE] */
                    {8'hbe,2'bx1} : dec_ma_enable = 1'b1;  /* XCH,A,[DE] */
                    {8'hbf,2'bx0} : dec_ma_enable = 1'b1;  /* XCH,A,[DE+byte] */
                    {8'hbf,2'bx1} : dec_ma_enable = 1'b1;  /* XCH,A,[DE+byte] */
                    {8'hbc,2'bx0} : dec_ma_enable = 1'b1;  /* XCH,A,[HL] */
                    {8'hbc,2'bx1} : dec_ma_enable = 1'b1;  /* XCH,A,[HL] */
                    {8'hbd,2'bx0} : dec_ma_enable = 1'b1;  /* XCH,A,[HL+byte] */
                    {8'hbd,2'bx1} : dec_ma_enable = 1'b1;  /* XCH,A,[HL+byte] */
                    {8'hd1,2'bxx} : dec_ma_enable = 1'b1;  /* AND,A,[HL+B] */
                    {8'he1,2'bxx} : dec_ma_enable = 1'b1;  /* OR,A,[HL+B] */
                    {8'hf1,2'bxx} : dec_ma_enable = 1'b1;  /* XOR,A,[HL+B] */
                    {8'h83,2'bxx} : dec_ma_enable = 1'b1;  /* ADD,A,[HL+C] */
                    {8'h93,2'bxx} : dec_ma_enable = 1'b1;  /* ADDC,A,[HL+C] */
                    {8'ha3,2'bxx} : dec_ma_enable = 1'b1;  /* SUB,A,[HL+C] */
                    {8'hb3,2'bxx} : dec_ma_enable = 1'b1;  /* SUBC,A,[HL+C] */
                    default : dec_ma_enable = 1'b0;
                endcase
            end else if(ID_stage0 == 8'h71) begin
                casex ({ID_stage1,stage_adr})  
                    {8'h04,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,saddr.0 */
                    {8'h14,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,saddr.1 */
                    {8'h24,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,saddr.2 */
                    {8'h34,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,saddr.3 */
                    {8'h44,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,saddr.4 */
                    {8'h54,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,saddr.5 */
                    {8'h64,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,saddr.6 */
                    {8'h74,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,saddr.7 */
                    {8'h0c,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,sfr.0 */
                    {8'h1c,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,sfr.1 */
                    {8'h2c,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,sfr.2 */
                    {8'h3c,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,sfr.3 */
                    {8'h4c,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,sfr.4 */
                    {8'h5c,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,sfr.5 */
                    {8'h6c,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,sfr.6 */
                    {8'h7c,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,sfr.7 */
                    {8'h84,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,[HL].0 */
                    {8'h94,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,[HL].1 */
                    {8'ha4,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,[HL].2 */
                    {8'hb4,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,[HL].3 */
                    {8'hc4,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,[HL].4 */
                    {8'hd4,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,[HL].5 */
                    {8'he4,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,[HL].6 */
                    {8'hf4,2'bxx} : dec_ma_enable = 1'b1;  /* MOV1,CY,[HL].7 */
                    {8'h01,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,saddr.0,CY */
                    {8'h01,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,saddr.0,CY */
                    {8'h11,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,saddr.1,CY */
                    {8'h11,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,saddr.1,CY */
                    {8'h21,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,saddr.2,CY */
                    {8'h21,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,saddr.2,CY */
                    {8'h31,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,saddr.3,CY */
                    {8'h31,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,saddr.3,CY */
                    {8'h41,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,saddr.4,CY */
                    {8'h41,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,saddr.4,CY */
                    {8'h51,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,saddr.5,CY */
                    {8'h51,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,saddr.5,CY */
                    {8'h61,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,saddr.6,CY */
                    {8'h61,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,saddr.6,CY */
                    {8'h71,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,saddr.7,CY */
                    {8'h71,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,saddr.7,CY */
                    {8'h09,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,sfr.0,CY */
                    {8'h09,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,sfr.0,CY */
                    {8'h19,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,sfr.1,CY */
                    {8'h19,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,sfr.1,CY */
                    {8'h29,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,sfr.2,CY */
                    {8'h29,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,sfr.2,CY */
                    {8'h39,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,sfr.3,CY */
                    {8'h39,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,sfr.3,CY */
                    {8'h49,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,sfr.4,CY */
                    {8'h49,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,sfr.4,CY */
                    {8'h59,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,sfr.5,CY */
                    {8'h59,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,sfr.5,CY */
                    {8'h69,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,sfr.6,CY */
                    {8'h69,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,sfr.6,CY */
                    {8'h79,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,sfr.7,CY */
                    {8'h79,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,sfr.7,CY */
                    {8'h81,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,[HL].0,CY */
                    {8'h81,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,[HL].0,CY */
                    {8'h91,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,[HL].1,CY */
                    {8'h91,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,[HL].1,CY */
                    {8'ha1,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,[HL].2,CY */
                    {8'ha1,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,[HL].2,CY */
                    {8'hb1,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,[HL].3,CY */
                    {8'hb1,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,[HL].3,CY */
                    {8'hc1,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,[HL].4,CY */
                    {8'hc1,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,[HL].4,CY */
                    {8'hd1,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,[HL].5,CY */
                    {8'hd1,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,[HL].5,CY */
                    {8'he1,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,[HL].6,CY */
                    {8'he1,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,[HL].6,CY */
                    {8'hf1,2'bx0} : dec_ma_enable = 1'b1;  /* MOV1,[HL].7,CY */
                    {8'hf1,2'bx1} : dec_ma_enable = 1'b1;  /* MOV1,[HL].7,CY */
                    {8'h05,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,saddr.0 */
                    {8'h15,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,saddr.1 */
                    {8'h25,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,saddr.2 */
                    {8'h35,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,saddr.3 */
                    {8'h45,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,saddr.4 */
                    {8'h55,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,saddr.5 */
                    {8'h65,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,saddr.6 */
                    {8'h75,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,saddr.7 */
                    {8'h0d,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,sfr.0 */
                    {8'h1d,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,sfr.1 */
                    {8'h2d,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,sfr.2 */
                    {8'h3d,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,sfr.3 */
                    {8'h4d,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,sfr.4 */
                    {8'h5d,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,sfr.5 */
                    {8'h6d,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,sfr.6 */
                    {8'h7d,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,sfr.7 */
                    {8'h85,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,[HL].0 */
                    {8'h95,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,[HL].1 */
                    {8'ha5,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,[HL].2 */
                    {8'hb5,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,[HL].3 */
                    {8'hc5,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,[HL].4 */
                    {8'hd5,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,[HL].5 */
                    {8'he5,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,[HL].6 */
                    {8'hf5,2'bxx} : dec_ma_enable = 1'b1;  /* AND1,CY,[HL].7 */
                    {8'h06,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,saddr.0 */
                    {8'h16,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,saddr.1 */
                    {8'h26,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,saddr.2 */
                    {8'h36,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,saddr.3 */
                    {8'h46,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,saddr.4 */
                    {8'h56,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,saddr.5 */
                    {8'h66,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,saddr.6 */
                    {8'h76,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,saddr.7 */
                    {8'h0e,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,sfr.0 */
                    {8'h1e,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,sfr.1 */
                    {8'h2e,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,sfr.2 */
                    {8'h3e,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,sfr.3 */
                    {8'h4e,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,sfr.4 */
                    {8'h5e,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,sfr.5 */
                    {8'h6e,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,sfr.6 */
                    {8'h7e,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,sfr.7 */
                    {8'h86,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,[HL].0 */
                    {8'h96,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,[HL].1 */
                    {8'ha6,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,[HL].2 */
                    {8'hb6,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,[HL].3 */
                    {8'hc6,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,[HL].4 */
                    {8'hd6,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,[HL].5 */
                    {8'he6,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,[HL].6 */
                    {8'hf6,2'bxx} : dec_ma_enable = 1'b1;  /* OR1,CY,[HL].7 */
                    {8'h07,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,saddr.0 */
                    {8'h17,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,saddr.1 */
                    {8'h27,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,saddr.2 */
                    {8'h37,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,saddr.3 */
                    {8'h47,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,saddr.4 */
                    {8'h57,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,saddr.5 */
                    {8'h67,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,saddr.6 */
                    {8'h77,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,saddr.7 */
                    {8'h0f,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,sfr.0 */
                    {8'h1f,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,sfr.1 */
                    {8'h2f,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,sfr.2 */
                    {8'h3f,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,sfr.3 */
                    {8'h4f,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,sfr.4 */
                    {8'h5f,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,sfr.5 */
                    {8'h6f,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,sfr.6 */
                    {8'h7f,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,sfr.7 */
                    {8'h87,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,[HL].0 */
                    {8'h97,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,[HL].1 */
                    {8'ha7,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,[HL].2 */
                    {8'hb7,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,[HL].3 */
                    {8'hc7,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,[HL].4 */
                    {8'hd7,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,[HL].5 */
                    {8'he7,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,[HL].6 */
                    {8'hf7,2'bxx} : dec_ma_enable = 1'b1;  /* XOR1,CY,[HL].7 */
                    {8'h02,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,saddr.0 */
                    {8'h02,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,saddr.0 */
                    {8'h12,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,saddr.1 */
                    {8'h12,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,saddr.1 */
                    {8'h22,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,saddr.2 */
                    {8'h22,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,saddr.2 */
                    {8'h32,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,saddr.3 */
                    {8'h32,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,saddr.3 */
                    {8'h42,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,saddr.4 */
                    {8'h42,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,saddr.4 */
                    {8'h52,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,saddr.5 */
                    {8'h52,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,saddr.5 */
                    {8'h62,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,saddr.6 */
                    {8'h62,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,saddr.6 */
                    {8'h72,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,saddr.7 */
                    {8'h72,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,saddr.7 */
                    {8'h0a,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,sfr.0 */
                    {8'h0a,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,sfr.0 */
                    {8'h1a,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,sfr.1 */
                    {8'h1a,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,sfr.1 */
                    {8'h2a,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,sfr.2 */
                    {8'h2a,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,sfr.2 */
                    {8'h3a,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,sfr.3 */
                    {8'h3a,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,sfr.3 */
                    {8'h4a,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,sfr.4 */
                    {8'h4a,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,sfr.4 */
                    {8'h5a,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,sfr.5 */
                    {8'h5a,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,sfr.5 */
                    {8'h6a,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,sfr.6 */
                    {8'h6a,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,sfr.6 */
                    {8'h7a,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,sfr.7 */
                    {8'h7a,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,sfr.7 */
                    {8'h00,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,!addr16.0 */
                    {8'h00,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,!addr16.0 */
                    {8'h10,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,!addr16.1 */
                    {8'h10,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,!addr16.1 */
                    {8'h20,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,!addr16.2 */
                    {8'h20,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,!addr16.2 */
                    {8'h30,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,!addr16.3 */
                    {8'h30,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,!addr16.3 */
                    {8'h40,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,!addr16.4 */
                    {8'h40,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,!addr16.4 */
                    {8'h50,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,!addr16.5 */
                    {8'h50,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,!addr16.5 */
                    {8'h60,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,!addr16.6 */
                    {8'h60,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,!addr16.6 */
                    {8'h70,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,!addr16.7 */
                    {8'h70,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,!addr16.7 */
                    {8'h82,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,[HL].0 */
                    {8'h82,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,[HL].0 */
                    {8'h92,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,[HL].1 */
                    {8'h92,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,[HL].1 */
                    {8'ha2,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,[HL].2 */
                    {8'ha2,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,[HL].2 */
                    {8'hb2,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,[HL].3 */
                    {8'hb2,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,[HL].3 */
                    {8'hc2,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,[HL].4 */
                    {8'hc2,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,[HL].4 */
                    {8'hd2,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,[HL].5 */
                    {8'hd2,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,[HL].5 */
                    {8'he2,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,[HL].6 */
                    {8'he2,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,[HL].6 */
                    {8'hf2,2'bx0} : dec_ma_enable = 1'b1;  /* SET1,,[HL].7 */
                    {8'hf2,2'bx1} : dec_ma_enable = 1'b1;  /* SET1,,[HL].7 */
                    {8'h03,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,saddr.0 */
                    {8'h03,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,saddr.0 */
                    {8'h13,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,saddr.1 */
                    {8'h13,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,saddr.1 */
                    {8'h23,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,saddr.2 */
                    {8'h23,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,saddr.2 */
                    {8'h33,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,saddr.3 */
                    {8'h33,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,saddr.3 */
                    {8'h43,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,saddr.4 */
                    {8'h43,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,saddr.4 */
                    {8'h53,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,saddr.5 */
                    {8'h53,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,saddr.5 */
                    {8'h63,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,saddr.6 */
                    {8'h63,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,saddr.6 */
                    {8'h73,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,saddr.7 */
                    {8'h73,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,saddr.7 */
                    {8'h0b,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,sfr.0 */
                    {8'h0b,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,sfr.0 */
                    {8'h1b,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,sfr.1 */
                    {8'h1b,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,sfr.1 */
                    {8'h2b,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,sfr.2 */
                    {8'h2b,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,sfr.2 */
                    {8'h3b,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,sfr.3 */
                    {8'h3b,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,sfr.3 */
                    {8'h4b,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,sfr.4 */
                    {8'h4b,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,sfr.4 */
                    {8'h5b,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,sfr.5 */
                    {8'h5b,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,sfr.5 */
                    {8'h6b,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,sfr.6 */
                    {8'h6b,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,sfr.6 */
                    {8'h7b,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,sfr.7 */
                    {8'h7b,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,sfr.7 */
                    {8'h08,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,!addr16.0 */
                    {8'h08,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,!addr16.0 */
                    {8'h18,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,!addr16.1 */
                    {8'h18,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,!addr16.1 */
                    {8'h28,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,!addr16.2 */
                    {8'h28,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,!addr16.2 */
                    {8'h38,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,!addr16.3 */
                    {8'h38,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,!addr16.3 */
                    {8'h48,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,!addr16.4 */
                    {8'h48,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,!addr16.4 */
                    {8'h58,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,!addr16.5 */
                    {8'h58,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,!addr16.5 */
                    {8'h68,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,!addr16.6 */
                    {8'h68,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,!addr16.6 */
                    {8'h78,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,!addr16.7 */
                    {8'h78,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,!addr16.7 */
                    {8'h83,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,[HL].0 */
                    {8'h83,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,[HL].0 */
                    {8'h93,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,[HL].1 */
                    {8'h93,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,[HL].1 */
                    {8'ha3,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,[HL].2 */
                    {8'ha3,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,[HL].2 */
                    {8'hb3,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,[HL].3 */
                    {8'hb3,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,[HL].3 */
                    {8'hc3,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,[HL].4 */
                    {8'hc3,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,[HL].4 */
                    {8'hd3,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,[HL].5 */
                    {8'hd3,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,[HL].5 */
                    {8'he3,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,[HL].6 */
                    {8'he3,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,[HL].6 */
                    {8'hf3,2'bx0} : dec_ma_enable = 1'b1;  /* CLR1,,[HL].7 */
                    {8'hf3,2'bx1} : dec_ma_enable = 1'b1;  /* CLR1,,[HL].7 */
                    default : dec_ma_enable = 1'b0;
                endcase
            end else if(ID_stage0 == 8'h31) begin
                casex ({ID_stage1,stage_adr})  
                    {8'h02,2'b00} : dec_ma_enable = 1'b1;  /* BT,saddr.0,$addr8 */
                    {8'h02,2'b01} : dec_ma_enable = 1'b1;  /* BT,saddr.0,$addr8 */
                    {8'h12,2'b00} : dec_ma_enable = 1'b1;  /* BT,saddr.1,$addr8 */
                    {8'h12,2'b01} : dec_ma_enable = 1'b1;  /* BT,saddr.1,$addr8 */
                    {8'h22,2'b00} : dec_ma_enable = 1'b1;  /* BT,saddr.2,$addr8 */
                    {8'h22,2'b01} : dec_ma_enable = 1'b1;  /* BT,saddr.2,$addr8 */
                    {8'h32,2'b00} : dec_ma_enable = 1'b1;  /* BT,saddr.3,$addr8 */
                    {8'h32,2'b01} : dec_ma_enable = 1'b1;  /* BT,saddr.3,$addr8 */
                    {8'h42,2'b00} : dec_ma_enable = 1'b1;  /* BT,saddr.4,$addr8 */
                    {8'h42,2'b01} : dec_ma_enable = 1'b1;  /* BT,saddr.4,$addr8 */
                    {8'h52,2'b00} : dec_ma_enable = 1'b1;  /* BT,saddr.5,$addr8 */
                    {8'h52,2'b01} : dec_ma_enable = 1'b1;  /* BT,saddr.5,$addr8 */
                    {8'h62,2'b00} : dec_ma_enable = 1'b1;  /* BT,saddr.6,$addr8 */
                    {8'h62,2'b01} : dec_ma_enable = 1'b1;  /* BT,saddr.6,$addr8 */
                    {8'h72,2'b00} : dec_ma_enable = 1'b1;  /* BT,saddr.7,$addr8 */
                    {8'h72,2'b01} : dec_ma_enable = 1'b1;  /* BT,saddr.7,$addr8 */
                    {8'h82,2'b00} : dec_ma_enable = 1'b1;  /* BT,sfr.0,$addr8 */
                    {8'h82,2'b01} : dec_ma_enable = 1'b1;  /* BT,sfr.0,$addr8 */
                    {8'h92,2'b00} : dec_ma_enable = 1'b1;  /* BT,sfr.1,$addr8 */
                    {8'h92,2'b01} : dec_ma_enable = 1'b1;  /* BT,sfr.1,$addr8 */
                    {8'ha2,2'b00} : dec_ma_enable = 1'b1;  /* BT,sfr.2,$addr8 */
                    {8'ha2,2'b01} : dec_ma_enable = 1'b1;  /* BT,sfr.2,$addr8 */
                    {8'hb2,2'b00} : dec_ma_enable = 1'b1;  /* BT,sfr.3,$addr8 */
                    {8'hb2,2'b01} : dec_ma_enable = 1'b1;  /* BT,sfr.3,$addr8 */
                    {8'hc2,2'b00} : dec_ma_enable = 1'b1;  /* BT,sfr.4,$addr8 */
                    {8'hc2,2'b01} : dec_ma_enable = 1'b1;  /* BT,sfr.4,$addr8 */
                    {8'hd2,2'b00} : dec_ma_enable = 1'b1;  /* BT,sfr.5,$addr8 */
                    {8'hd2,2'b01} : dec_ma_enable = 1'b1;  /* BT,sfr.5,$addr8 */
                    {8'he2,2'b00} : dec_ma_enable = 1'b1;  /* BT,sfr.6,$addr8 */
                    {8'he2,2'b01} : dec_ma_enable = 1'b1;  /* BT,sfr.6,$addr8 */
                    {8'hf2,2'b00} : dec_ma_enable = 1'b1;  /* BT,sfr.7,$addr8 */
                    {8'hf2,2'b01} : dec_ma_enable = 1'b1;  /* BT,sfr.7,$addr8 */
                    {8'h83,2'b00} : dec_ma_enable = 1'b1;  /* BT,[HL].0,$addr8 */
                    {8'h83,2'b01} : dec_ma_enable = 1'b1;  /* BT,[HL].0,$addr8 */
                    {8'h93,2'b00} : dec_ma_enable = 1'b1;  /* BT,[HL].1,$addr8 */
                    {8'h93,2'b01} : dec_ma_enable = 1'b1;  /* BT,[HL].1,$addr8 */
                    {8'ha3,2'b00} : dec_ma_enable = 1'b1;  /* BT,[HL].2,$addr8 */
                    {8'ha3,2'b01} : dec_ma_enable = 1'b1;  /* BT,[HL].2,$addr8 */
                    {8'hb3,2'b00} : dec_ma_enable = 1'b1;  /* BT,[HL].3,$addr8 */
                    {8'hb3,2'b01} : dec_ma_enable = 1'b1;  /* BT,[HL].3,$addr8 */
                    {8'hc3,2'b00} : dec_ma_enable = 1'b1;  /* BT,[HL].4,$addr8 */
                    {8'hc3,2'b01} : dec_ma_enable = 1'b1;  /* BT,[HL].4,$addr8 */
                    {8'hd3,2'b00} : dec_ma_enable = 1'b1;  /* BT,[HL].5,$addr8 */
                    {8'hd3,2'b01} : dec_ma_enable = 1'b1;  /* BT,[HL].5,$addr8 */
                    {8'he3,2'b00} : dec_ma_enable = 1'b1;  /* BT,[HL].6,$addr8 */
                    {8'he3,2'b01} : dec_ma_enable = 1'b1;  /* BT,[HL].6,$addr8 */
                    {8'hf3,2'b00} : dec_ma_enable = 1'b1;  /* BT,[HL].7,$addr8 */
                    {8'hf3,2'b01} : dec_ma_enable = 1'b1;  /* BT,[HL].7,$addr8 */
                    {8'h04,2'b00} : dec_ma_enable = 1'b1;  /* BF,saddr.0,$addr8 */
                    {8'h04,2'b01} : dec_ma_enable = 1'b1;  /* BF,saddr.0,$addr8 */
                    {8'h14,2'b00} : dec_ma_enable = 1'b1;  /* BF,saddr.1,$addr8 */
                    {8'h14,2'b01} : dec_ma_enable = 1'b1;  /* BF,saddr.1,$addr8 */
                    {8'h24,2'b00} : dec_ma_enable = 1'b1;  /* BF,saddr.2,$addr8 */
                    {8'h24,2'b01} : dec_ma_enable = 1'b1;  /* BF,saddr.2,$addr8 */
                    {8'h34,2'b00} : dec_ma_enable = 1'b1;  /* BF,saddr.3,$addr8 */
                    {8'h34,2'b01} : dec_ma_enable = 1'b1;  /* BF,saddr.3,$addr8 */
                    {8'h44,2'b00} : dec_ma_enable = 1'b1;  /* BF,saddr.4,$addr8 */
                    {8'h44,2'b01} : dec_ma_enable = 1'b1;  /* BF,saddr.4,$addr8 */
                    {8'h54,2'b00} : dec_ma_enable = 1'b1;  /* BF,saddr.5,$addr8 */
                    {8'h54,2'b01} : dec_ma_enable = 1'b1;  /* BF,saddr.5,$addr8 */
                    {8'h64,2'b00} : dec_ma_enable = 1'b1;  /* BF,saddr.6,$addr8 */
                    {8'h64,2'b01} : dec_ma_enable = 1'b1;  /* BF,saddr.6,$addr8 */
                    {8'h74,2'b00} : dec_ma_enable = 1'b1;  /* BF,saddr.7,$addr8 */
                    {8'h74,2'b01} : dec_ma_enable = 1'b1;  /* BF,saddr.7,$addr8 */
                    {8'h84,2'b00} : dec_ma_enable = 1'b1;  /* BF,sfr.0,$addr8 */
                    {8'h84,2'b01} : dec_ma_enable = 1'b1;  /* BF,sfr.0,$addr8 */
                    {8'h94,2'b00} : dec_ma_enable = 1'b1;  /* BF,sfr.1,$addr8 */
                    {8'h94,2'b01} : dec_ma_enable = 1'b1;  /* BF,sfr.1,$addr8 */
                    {8'ha4,2'b00} : dec_ma_enable = 1'b1;  /* BF,sfr.2,$addr8 */
                    {8'ha4,2'b01} : dec_ma_enable = 1'b1;  /* BF,sfr.2,$addr8 */
                    {8'hb4,2'b00} : dec_ma_enable = 1'b1;  /* BF,sfr.3,$addr8 */
                    {8'hb4,2'b01} : dec_ma_enable = 1'b1;  /* BF,sfr.3,$addr8 */
                    {8'hc4,2'b00} : dec_ma_enable = 1'b1;  /* BF,sfr.4,$addr8 */
                    {8'hc4,2'b01} : dec_ma_enable = 1'b1;  /* BF,sfr.4,$addr8 */
                    {8'hd4,2'b00} : dec_ma_enable = 1'b1;  /* BF,sfr.5,$addr8 */
                    {8'hd4,2'b01} : dec_ma_enable = 1'b1;  /* BF,sfr.5,$addr8 */
                    {8'he4,2'b00} : dec_ma_enable = 1'b1;  /* BF,sfr.6,$addr8 */
                    {8'he4,2'b01} : dec_ma_enable = 1'b1;  /* BF,sfr.6,$addr8 */
                    {8'hf4,2'b00} : dec_ma_enable = 1'b1;  /* BF,sfr.7,$addr8 */
                    {8'hf4,2'b01} : dec_ma_enable = 1'b1;  /* BF,sfr.7,$addr8 */
                    {8'h85,2'b00} : dec_ma_enable = 1'b1;  /* BF,[HL].0,$addr8 */
                    {8'h85,2'b01} : dec_ma_enable = 1'b1;  /* BF,[HL].0,$addr8 */
                    {8'h95,2'b00} : dec_ma_enable = 1'b1;  /* BF,[HL].1,$addr8 */
                    {8'h95,2'b01} : dec_ma_enable = 1'b1;  /* BF,[HL].1,$addr8 */
                    {8'ha5,2'b00} : dec_ma_enable = 1'b1;  /* BF,[HL].2,$addr8 */
                    {8'ha5,2'b01} : dec_ma_enable = 1'b1;  /* BF,[HL].2,$addr8 */
                    {8'hb5,2'b00} : dec_ma_enable = 1'b1;  /* BF,[HL].3,$addr8 */
                    {8'hb5,2'b01} : dec_ma_enable = 1'b1;  /* BF,[HL].3,$addr8 */
                    {8'hc5,2'b00} : dec_ma_enable = 1'b1;  /* BF,[HL].4,$addr8 */
                    {8'hc5,2'b01} : dec_ma_enable = 1'b1;  /* BF,[HL].4,$addr8 */
                    {8'hd5,2'b00} : dec_ma_enable = 1'b1;  /* BF,[HL].5,$addr8 */
                    {8'hd5,2'b01} : dec_ma_enable = 1'b1;  /* BF,[HL].5,$addr8 */
                    {8'he5,2'b00} : dec_ma_enable = 1'b1;  /* BF,[HL].6,$addr8 */
                    {8'he5,2'b01} : dec_ma_enable = 1'b1;  /* BF,[HL].6,$addr8 */
                    {8'hf5,2'b00} : dec_ma_enable = 1'b1;  /* BF,[HL].7,$addr8 */
                    {8'hf5,2'b01} : dec_ma_enable = 1'b1;  /* BF,[HL].7,$addr8 */
                    {8'h00,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.0,$addr8 */
                    {8'h00,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.0,$addr8 */
                    {8'h00,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.0,$addr8 */
                    {8'h10,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.1,$addr8 */
                    {8'h10,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.1,$addr8 */
                    {8'h10,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.1,$addr8 */
                    {8'h20,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.2,$addr8 */
                    {8'h20,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.2,$addr8 */
                    {8'h20,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.2,$addr8 */
                    {8'h30,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.3,$addr8 */
                    {8'h30,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.3,$addr8 */
                    {8'h30,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.3,$addr8 */
                    {8'h40,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.4,$addr8 */
                    {8'h40,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.4,$addr8 */
                    {8'h40,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.4,$addr8 */
                    {8'h50,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.5,$addr8 */
                    {8'h50,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.5,$addr8 */
                    {8'h50,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.5,$addr8 */
                    {8'h60,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.6,$addr8 */
                    {8'h60,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.6,$addr8 */
                    {8'h60,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.6,$addr8 */
                    {8'h70,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.7,$addr8 */
                    {8'h70,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.7,$addr8 */
                    {8'h70,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,saddr.7,$addr8 */
                    {8'h80,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.0,$addr8 */
                    {8'h80,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.0,$addr8 */
                    {8'h80,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.0,$addr8 */
                    {8'h90,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.1,$addr8 */
                    {8'h90,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.1,$addr8 */
                    {8'h90,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.1,$addr8 */
                    {8'ha0,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.2,$addr8 */
                    {8'ha0,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.2,$addr8 */
                    {8'ha0,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.2,$addr8 */
                    {8'hb0,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.3,$addr8 */
                    {8'hb0,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.3,$addr8 */
                    {8'hb0,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.3,$addr8 */
                    {8'hc0,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.4,$addr8 */
                    {8'hc0,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.4,$addr8 */
                    {8'hc0,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.4,$addr8 */
                    {8'hd0,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.5,$addr8 */
                    {8'hd0,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.5,$addr8 */
                    {8'hd0,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.5,$addr8 */
                    {8'he0,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.6,$addr8 */
                    {8'he0,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.6,$addr8 */
                    {8'he0,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.6,$addr8 */
                    {8'hf0,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.7,$addr8 */
                    {8'hf0,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.7,$addr8 */
                    {8'hf0,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,sfr.7,$addr8 */
                    {8'h81,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].0,$addr8 */
                    {8'h81,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].0,$addr8 */
                    {8'h81,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].0,$addr8 */
                    {8'h91,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].1,$addr8 */
                    {8'h91,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].1,$addr8 */
                    {8'h91,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].1,$addr8 */
                    {8'ha1,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].2,$addr8 */
                    {8'ha1,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].2,$addr8 */
                    {8'ha1,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].2,$addr8 */
                    {8'hb1,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].3,$addr8 */
                    {8'hb1,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].3,$addr8 */
                    {8'hb1,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].3,$addr8 */
                    {8'hc1,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].4,$addr8 */
                    {8'hc1,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].4,$addr8 */
                    {8'hc1,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].4,$addr8 */
                    {8'hd1,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].5,$addr8 */
                    {8'hd1,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].5,$addr8 */
                    {8'hd1,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].5,$addr8 */
                    {8'he1,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].6,$addr8 */
                    {8'he1,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].6,$addr8 */
                    {8'he1,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].6,$addr8 */
                    {8'hf1,2'b00} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].7,$addr8 */
                    {8'hf1,2'b01} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].7,$addr8 */
                    {8'hf1,2'b10} : dec_ma_enable = 1'b1;  /* BTCLR,[HL].7,$addr8 */
                    default : dec_ma_enable = 1'b0;
                endcase
            end else begin
                casex ({ID_stage0,stage_adr})  
                    {8'hcd,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,saddr,#byte */
                    {8'hce,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,sfr,#byte */
                    {8'hcf,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,!addr16,#byte */
                    {8'hca,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,[DE+byte],#byte */
                    {8'hcc,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,[HL+byte],#byte */
                    {8'h8d,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,A,saddr */
                    {8'h9d,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,saddr,A */
                    {8'h8e,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,A,sfr */
                    {8'h9e,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,sfr,A */
                    {8'h8f,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,A,!addr16 */
                    {8'h9f,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,!addr16,A */
                    {8'h89,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,A,[DE] */
                    {8'h99,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,[DE],A */
                    {8'h8a,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,A,[DE+byte] */
                    {8'h9a,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,[DE+byte],A */
                    {8'h8b,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,A,[HL] */
                    {8'h9b,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,[HL],A */
                    {8'h8c,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,A,[HL+byte] */
                    {8'h9c,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,[HL+byte],A */
                    {8'h19,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,word[B],#byte */
                    {8'h09,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,A,word[B] */
                    {8'h18,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,word[B],A */
                    {8'h38,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,word[C],#byte */
                    {8'h29,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,A,word[C] */
                    {8'h28,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,word[C],A */
                    {8'h39,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,word[BC],#byte */
                    {8'h49,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,A,word[BC] */
                    {8'h48,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,word[BC],A */
                    {8'hc8,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,[SP+byte],#byte */
                    {8'h88,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,A,[SP+byte] */
                    {8'h98,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,[SP+byte],A */
                    {8'he8,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,B,saddr */
                    {8'he9,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,B,!addr16 */
                    {8'hf8,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,C,saddr */
                    {8'hf9,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,C,!addr16 */
                    {8'hd8,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,X,saddr */
                    {8'hd9,2'bxx} : dec_ma_enable = 1'b1;  /* MOV,X,!addr16 */
                    {8'he4,2'bxx} : dec_ma_enable = 1'b1;  /* ONEB,,saddr */
                    {8'he5,2'bxx} : dec_ma_enable = 1'b1;  /* ONEB,,!addr16 */
                    {8'hf4,2'bxx} : dec_ma_enable = 1'b1;  /* CLRB,,saddr */
                    {8'hf5,2'bxx} : dec_ma_enable = 1'b1;  /* CLRB,,!addr16 */
                    {8'hc9,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,saddrp,#word */
                    {8'hcb,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,sfrp,#word */
                    {8'had,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,AX,saddrp */
                    {8'hbd,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,saddrp,AX */
                    {8'hae,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,AX,sfrp */
                    {8'hbe,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,sfrp,AX */
                    {8'haf,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,AX,!addr16 */
                    {8'hbf,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,!addr16,AX */
                    {8'ha9,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,AX,[DE] */
                    {8'haa,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,AX,[DE+byte] */
                    {8'hb9,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,[DE],AX */
                    {8'hba,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,[DE+byte],AX */
                    {8'hab,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,AX,[HL] */
                    {8'hac,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,AX,[HL+byte] */
                    {8'hbb,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,[HL],AX */
                    {8'hbc,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,[HL+byte],AX */
                    {8'h59,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,AX,word[B] */
                    {8'h58,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,word[B],AX */
                    {8'h69,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,AX,word[C] */
                    {8'h68,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,word[C],AX */
                    {8'h79,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,AX,word[BC] */
                    {8'h78,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,word[BC],AX */
                    {8'ha8,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,AX,[SP+byte] */
                    {8'hb8,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,[SP+byte],AX */
                    {8'hda,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,BC,saddrp */
                    {8'hdb,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,BC,!addr16 */
                    {8'hea,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,DE,saddrp */
                    {8'heb,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,DE,!addr16 */
                    {8'hfa,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,HL,saddrp */
                    {8'hfb,2'bxx} : dec_ma_enable = 1'b1;  /* MOVW,HL,!addr16 */
                    {8'h0a,2'bx0} : dec_ma_enable = 1'b1;  /* ADD,saddr,#byte */
                    {8'h0a,2'bx1} : dec_ma_enable = 1'b1;  /* ADD,saddr,#byte */
                    {8'h0b,2'bxx} : dec_ma_enable = 1'b1;  /* ADD,A,saddr */
                    {8'h0f,2'bxx} : dec_ma_enable = 1'b1;  /* ADD,A,!addr16 */
                    {8'h0d,2'bxx} : dec_ma_enable = 1'b1;  /* ADD,A,[HL] */
                    {8'h0e,2'bxx} : dec_ma_enable = 1'b1;  /* ADD,A,[HL+byte] */
                    {8'h1a,2'bx0} : dec_ma_enable = 1'b1;  /* ADDC,saddr,#byte */
                    {8'h1a,2'bx1} : dec_ma_enable = 1'b1;  /* ADDC,saddr,#byte */
                    {8'h1b,2'bxx} : dec_ma_enable = 1'b1;  /* ADDC,A,saddr */
                    {8'h1f,2'bxx} : dec_ma_enable = 1'b1;  /* ADDC,A,!addr16 */
                    {8'h1d,2'bxx} : dec_ma_enable = 1'b1;  /* ADDC,A,[HL] */
                    {8'h1e,2'bxx} : dec_ma_enable = 1'b1;  /* ADDC,A,[HL+byte] */
                    {8'h2a,2'bx0} : dec_ma_enable = 1'b1;  /* SUB,saddr,#byte */
                    {8'h2a,2'bx1} : dec_ma_enable = 1'b1;  /* SUB,saddr,#byte */
                    {8'h2b,2'bxx} : dec_ma_enable = 1'b1;  /* SUB,A,saddr */
                    {8'h2f,2'bxx} : dec_ma_enable = 1'b1;  /* SUB,A,!addr16 */
                    {8'h2d,2'bxx} : dec_ma_enable = 1'b1;  /* SUB,A,[HL] */
                    {8'h2e,2'bxx} : dec_ma_enable = 1'b1;  /* SUB,A,[HL+byte] */
                    {8'h3a,2'bx0} : dec_ma_enable = 1'b1;  /* SUBC,saddr,#byte */
                    {8'h3a,2'bx1} : dec_ma_enable = 1'b1;  /* SUBC,saddr,#byte */
                    {8'h3b,2'bxx} : dec_ma_enable = 1'b1;  /* SUBC,A,saddr */
                    {8'h3f,2'bxx} : dec_ma_enable = 1'b1;  /* SUBC,A,!addr16 */
                    {8'h3d,2'bxx} : dec_ma_enable = 1'b1;  /* SUBC,A,[HL] */
                    {8'h3e,2'bxx} : dec_ma_enable = 1'b1;  /* SUBC,A,[HL+byte] */
                    {8'h5a,2'bx0} : dec_ma_enable = 1'b1;  /* AND,saddr,#byte */
                    {8'h5a,2'bx1} : dec_ma_enable = 1'b1;  /* AND,saddr,#byte */
                    {8'h5b,2'bxx} : dec_ma_enable = 1'b1;  /* AND,A,saddr */
                    {8'h5f,2'bxx} : dec_ma_enable = 1'b1;  /* AND,A,!addr16 */
                    {8'h5d,2'bxx} : dec_ma_enable = 1'b1;  /* AND,A,[HL] */
                    {8'h5e,2'bxx} : dec_ma_enable = 1'b1;  /* AND,A,[HL+byte] */
                    {8'h6a,2'bx0} : dec_ma_enable = 1'b1;  /* OR,saddr,#byte */
                    {8'h6a,2'bx1} : dec_ma_enable = 1'b1;  /* OR,saddr,#byte */
                    {8'h6b,2'bxx} : dec_ma_enable = 1'b1;  /* OR,A,saddr */
                    {8'h6f,2'bxx} : dec_ma_enable = 1'b1;  /* OR,A,!addr16 */
                    {8'h6d,2'bxx} : dec_ma_enable = 1'b1;  /* OR,A,[HL] */
                    {8'h6e,2'bxx} : dec_ma_enable = 1'b1;  /* OR,A,[HL+byte] */
                    {8'h7a,2'bx0} : dec_ma_enable = 1'b1;  /* XOR,saddr,#byte */
                    {8'h7a,2'bx1} : dec_ma_enable = 1'b1;  /* XOR,saddr,#byte */
                    {8'h7b,2'bxx} : dec_ma_enable = 1'b1;  /* XOR,A,saddr */
                    {8'h7f,2'bxx} : dec_ma_enable = 1'b1;  /* XOR,A,!addr16 */
                    {8'h7d,2'bxx} : dec_ma_enable = 1'b1;  /* XOR,A,[HL] */
                    {8'h7e,2'bxx} : dec_ma_enable = 1'b1;  /* XOR,A,[HL+byte] */
                    {8'h4a,2'bxx} : dec_ma_enable = 1'b1;  /* CMP,saddr,#byte */
                    {8'h40,2'bxx} : dec_ma_enable = 1'b1;  /* CMP,!addr16,#byte */
                    {8'h4b,2'bxx} : dec_ma_enable = 1'b1;  /* CMP,A,saddr */
                    {8'h4f,2'bxx} : dec_ma_enable = 1'b1;  /* CMP,A,!addr16 */
                    {8'h4d,2'bxx} : dec_ma_enable = 1'b1;  /* CMP,A,[HL] */
                    {8'h4e,2'bxx} : dec_ma_enable = 1'b1;  /* CMP,A,[HL+byte] */
                    {8'hd4,2'bxx} : dec_ma_enable = 1'b1;  /* CMP0,,saddr */
                    {8'hd5,2'bxx} : dec_ma_enable = 1'b1;  /* CMP0,,!addr16 */
                    {8'h06,2'bxx} : dec_ma_enable = 1'b1;  /* ADDW,AX,saddrp */
                    {8'h02,2'bxx} : dec_ma_enable = 1'b1;  /* ADDW,AX,!addr16 */
                    {8'h26,2'bxx} : dec_ma_enable = 1'b1;  /* SUBW,AX,saddrp */
                    {8'h22,2'bxx} : dec_ma_enable = 1'b1;  /* SUBW,AX,!addr16 */
                    {8'h46,2'bxx} : dec_ma_enable = 1'b1;  /* CMPW,AX,saddrp */
                    {8'h42,2'bxx} : dec_ma_enable = 1'b1;  /* CMPW,AX,!addr16 */
                    {8'ha4,2'bx0} : dec_ma_enable = 1'b1;  /* INC,,saddr */
                    {8'ha4,2'bx1} : dec_ma_enable = 1'b1;  /* INC,,saddr */
                    {8'ha0,2'bx0} : dec_ma_enable = 1'b1;  /* INC,,!addr16 */
                    {8'ha0,2'bx1} : dec_ma_enable = 1'b1;  /* INC,,!addr16 */
                    {8'hb4,2'bx0} : dec_ma_enable = 1'b1;  /* DEC,,saddr */
                    {8'hb4,2'bx1} : dec_ma_enable = 1'b1;  /* DEC,,saddr */
                    {8'hb0,2'bx0} : dec_ma_enable = 1'b1;  /* DEC,,!addr16 */
                    {8'hb0,2'bx1} : dec_ma_enable = 1'b1;  /* DEC,,!addr16 */
                    {8'ha6,2'bx0} : dec_ma_enable = 1'b1;  /* INCW,,saddrp */
                    {8'ha6,2'bx1} : dec_ma_enable = 1'b1;  /* INCW,,saddrp */
                    {8'ha2,2'bx0} : dec_ma_enable = 1'b1;  /* INCW,,!addr16 */
                    {8'ha2,2'bx1} : dec_ma_enable = 1'b1;  /* INCW,,!addr16 */
                    {8'hb6,2'bx0} : dec_ma_enable = 1'b1;  /* DECW,,saddrp */
                    {8'hb6,2'bx1} : dec_ma_enable = 1'b1;  /* DECW,,saddrp */
                    {8'hb2,2'bx0} : dec_ma_enable = 1'b1;  /* DECW,,!addr16 */
                    {8'hb2,2'bx1} : dec_ma_enable = 1'b1;  /* DECW,,!addr16 */
                    {8'hfe,2'bx0} : dec_ma_enable = 1'b1;  /* CALL,,$!addr16 */
                    {8'hfe,2'bx1} : dec_ma_enable = 1'b1;  /* CALL,,$!addr16 */
                    {8'hfd,2'bx0} : dec_ma_enable = 1'b1;  /* CALL,,!addr16 */
                    {8'hfd,2'bx1} : dec_ma_enable = 1'b1;  /* CALL,,!addr16 */
                    {8'hfc,2'bx0} : dec_ma_enable = 1'b1;  /* CALL,,!!addr20 */
                    {8'hfc,2'bx1} : dec_ma_enable = 1'b1;  /* CALL,,!!addr20 */
                    {8'hd7,2'b00} : dec_ma_enable = 1'b1;  /* RET,, */
                    {8'hd7,2'b01} : dec_ma_enable = 1'b1;  /* RET,, */
                    {8'hc1,2'bxx} : dec_ma_enable = 1'b1;  /* PUSH,,AX */
                    {8'hc3,2'bxx} : dec_ma_enable = 1'b1;  /* PUSH,,BC */
                    {8'hc5,2'bxx} : dec_ma_enable = 1'b1;  /* PUSH,,DE */
                    {8'hc7,2'bxx} : dec_ma_enable = 1'b1;  /* PUSH,,HL */
                    {8'hc0,2'bxx} : dec_ma_enable = 1'b1;  /* POP,,AX */
                    {8'hc2,2'bxx} : dec_ma_enable = 1'b1;  /* POP,,BC */
                    {8'hc4,2'bxx} : dec_ma_enable = 1'b1;  /* POP,,DE */
                    {8'hc6,2'bxx} : dec_ma_enable = 1'b1;  /* POP,,HL */
                    {8'hff,2'bx0} : dec_ma_enable = 1'b1;  /* SOFT,,BREAK */
                    {8'hff,2'bx1} : dec_ma_enable = 1'b1;  /* SOFT,,BREAK */
                    default : dec_ma_enable = 1'b0;
                endcase
            end
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ma_data_sp;
    reg    dec_ma_data_sp;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(decout_mask == 1'b1) begin
//            dec_ma_data_sp = 1'b0;
//        end else if(rstvec == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1) begin
            dec_ma_data_sp = 1'b0;
        end else if(ivack == 1'b1) begin
            casex ({stage_adr})  
                {2'b00} : dec_ma_data_sp = 1'b1;  /* Interrupt */
                {2'b01} : dec_ma_data_sp = 1'b1;  /* Interrupt */
                default : dec_ma_data_sp = 1'b0;
            endcase
        end else if(skpack == 1'b1) begin
            dec_ma_data_sp = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hca,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALL,,AX */
                {8'h61,8'hca,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALL,,AX */
                {8'h61,8'hda,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALL,,BC */
                {8'h61,8'hda,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALL,,BC */
                {8'h61,8'hea,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALL,,DE */
                {8'h61,8'hea,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALL,,DE */
                {8'h61,8'hfa,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALL,,HL */
                {8'h61,8'hfa,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALL,,HL */
                {8'hfe,8'hxx,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALL,,$!addr16 */
                {8'hfe,8'hxx,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALL,,$!addr16 */
                {8'hfd,8'hxx,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALL,,!addr16 */
                {8'hfd,8'hxx,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALL,,!addr16 */
                {8'hfc,8'hxx,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALL,,!!addr20 */
                {8'hfc,8'hxx,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALL,,!!addr20 */
                {8'h61,8'h84,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[0080h] */
                {8'h61,8'h84,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[0080h] */
                {8'h61,8'h94,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[0082h] */
                {8'h61,8'h94,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[0082h] */
                {8'h61,8'ha4,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[0084h] */
                {8'h61,8'ha4,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[0084h] */
                {8'h61,8'hb4,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[0086h] */
                {8'h61,8'hb4,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[0086h] */
                {8'h61,8'hc4,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[0088h] */
                {8'h61,8'hc4,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[0088h] */
                {8'h61,8'hd4,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[008Ah] */
                {8'h61,8'hd4,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[008Ah] */
                {8'h61,8'he4,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[008Ch] */
                {8'h61,8'he4,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[008Ch] */
                {8'h61,8'hf4,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[008Eh] */
                {8'h61,8'hf4,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[008Eh] */
                {8'h61,8'h85,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[0090h] */
                {8'h61,8'h85,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[0090h] */
                {8'h61,8'h95,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[0092h] */
                {8'h61,8'h95,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[0092h] */
                {8'h61,8'ha5,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[0094h] */
                {8'h61,8'ha5,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[0094h] */
                {8'h61,8'hb5,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[0096h] */
                {8'h61,8'hb5,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[0096h] */
                {8'h61,8'hc5,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[0098h] */
                {8'h61,8'hc5,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[0098h] */
                {8'h61,8'hd5,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[009Ah] */
                {8'h61,8'hd5,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[009Ah] */
                {8'h61,8'he5,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[009Ch] */
                {8'h61,8'he5,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[009Ch] */
                {8'h61,8'hf5,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[009Eh] */
                {8'h61,8'hf5,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[009Eh] */
                {8'h61,8'h86,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00A0h] */
                {8'h61,8'h86,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00A0h] */
                {8'h61,8'h96,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00A2h] */
                {8'h61,8'h96,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00A2h] */
                {8'h61,8'ha6,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00A4h] */
                {8'h61,8'ha6,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00A4h] */
                {8'h61,8'hb6,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00A6h] */
                {8'h61,8'hb6,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00A6h] */
                {8'h61,8'hc6,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00A8h] */
                {8'h61,8'hc6,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00A8h] */
                {8'h61,8'hd6,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00AAh] */
                {8'h61,8'hd6,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00AAh] */
                {8'h61,8'he6,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00ACh] */
                {8'h61,8'he6,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00ACh] */
                {8'h61,8'hf6,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00AEh] */
                {8'h61,8'hf6,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00AEh] */
                {8'h61,8'h87,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00B0h] */
                {8'h61,8'h87,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00B0h] */
                {8'h61,8'h97,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00B2h] */
                {8'h61,8'h97,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00B2h] */
                {8'h61,8'ha7,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00B4h] */
                {8'h61,8'ha7,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00B4h] */
                {8'h61,8'hb7,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00B6h] */
                {8'h61,8'hb7,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00B6h] */
                {8'h61,8'hc7,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00B8h] */
                {8'h61,8'hc7,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00B8h] */
                {8'h61,8'hd7,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00BAh] */
                {8'h61,8'hd7,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00BAh] */
                {8'h61,8'he7,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00BCh] */
                {8'h61,8'he7,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00BCh] */
                {8'h61,8'hf7,2'bx0} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00BEh] */
                {8'h61,8'hf7,2'bx1} : dec_ma_data_sp = 1'b1;  /* CALLT,,[00BEh] */
                {8'h61,8'hcc,2'bx0} : dec_ma_data_sp = 1'b1;  /* BRK,, */
                {8'h61,8'hcc,2'bx1} : dec_ma_data_sp = 1'b1;  /* BRK,, */
                {8'hd7,8'hxx,2'b00} : dec_ma_data_sp = 1'b1;  /* RET,, */
                {8'hd7,8'hxx,2'b01} : dec_ma_data_sp = 1'b1;  /* RET,, */
                {8'h61,8'hec,2'b00} : dec_ma_data_sp = 1'b1;  /* RETB,, */
                {8'h61,8'hec,2'b01} : dec_ma_data_sp = 1'b1;  /* RETB,, */
                {8'h61,8'hfc,2'b00} : dec_ma_data_sp = 1'b1;  /* RETI,, */
                {8'h61,8'hfc,2'b01} : dec_ma_data_sp = 1'b1;  /* RETI,, */
                {8'h61,8'hdd,2'bxx} : dec_ma_data_sp = 1'b1;  /* PUSH,,PSW */
                {8'hc1,8'hxx,2'bxx} : dec_ma_data_sp = 1'b1;  /* PUSH,,AX */
                {8'hc3,8'hxx,2'bxx} : dec_ma_data_sp = 1'b1;  /* PUSH,,BC */
                {8'hc5,8'hxx,2'bxx} : dec_ma_data_sp = 1'b1;  /* PUSH,,DE */
                {8'hc7,8'hxx,2'bxx} : dec_ma_data_sp = 1'b1;  /* PUSH,,HL */
                {8'h61,8'hcd,2'bxx} : dec_ma_data_sp = 1'b1;  /* POP,,PSW */
                {8'hc0,8'hxx,2'bxx} : dec_ma_data_sp = 1'b1;  /* POP,,AX */
                {8'hc2,8'hxx,2'bxx} : dec_ma_data_sp = 1'b1;  /* POP,,BC */
                {8'hc4,8'hxx,2'bxx} : dec_ma_data_sp = 1'b1;  /* POP,,DE */
                {8'hc6,8'hxx,2'bxx} : dec_ma_data_sp = 1'b1;  /* POP,,HL */
                {8'hff,8'hxx,2'bx0} : dec_ma_data_sp = 1'b1;  /* SOFT,,BREAK */
                {8'hff,8'hxx,2'bx1} : dec_ma_data_sp = 1'b1;  /* SOFT,,BREAK */
                {8'h61,8'ha1,2'bx0} : dec_ma_data_sp = 1'b1;  /* SOFT2,,BREAK */
                {8'h61,8'ha1,2'bx1} : dec_ma_data_sp = 1'b1;  /* SOFT2,,BREAK */
                {8'h61,8'hb1,2'bx0} : dec_ma_data_sp = 1'b1;  /* SOFT3,,BREAK */
                {8'h61,8'hb1,2'bx1} : dec_ma_data_sp = 1'b1;  /* SOFT3,,BREAK */
                {8'h61,8'hc1,2'bx0} : dec_ma_data_sp = 1'b1;  /* SOFT4,,BREAK */
                {8'h61,8'hc1,2'bx1} : dec_ma_data_sp = 1'b1;  /* SOFT4,,BREAK */
                default : dec_ma_data_sp = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ma_data_saddr_op1;
    reg    dec_ma_data_saddr_op1;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_ma_data_saddr_op1 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'hcd,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* MOV,saddr,#byte */
                {8'h8d,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* MOV,A,saddr */
                {8'h9d,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* MOV,saddr,A */
                {8'he8,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* MOV,B,saddr */
                {8'hf8,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* MOV,C,saddr */
                {8'hd8,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* MOV,X,saddr */
                {8'he4,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* ONEB,,saddr */
                {8'hf4,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* CLRB,,saddr */
                {8'hc9,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* MOVW,saddrp,#word */
                {8'had,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* MOVW,AX,saddrp */
                {8'hbd,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* MOVW,saddrp,AX */
                {8'hda,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* MOVW,BC,saddrp */
                {8'hea,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* MOVW,DE,saddrp */
                {8'hfa,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* MOVW,HL,saddrp */
                {8'h0a,8'hxx,2'bx0} : dec_ma_data_saddr_op1 = 1'b1;  /* ADD,saddr,#byte */
                {8'h0a,8'hxx,2'bx1} : dec_ma_data_saddr_op1 = 1'b1;  /* ADD,saddr,#byte */
                {8'h0b,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* ADD,A,saddr */
                {8'h1a,8'hxx,2'bx0} : dec_ma_data_saddr_op1 = 1'b1;  /* ADDC,saddr,#byte */
                {8'h1a,8'hxx,2'bx1} : dec_ma_data_saddr_op1 = 1'b1;  /* ADDC,saddr,#byte */
                {8'h1b,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* ADDC,A,saddr */
                {8'h2a,8'hxx,2'bx0} : dec_ma_data_saddr_op1 = 1'b1;  /* SUB,saddr,#byte */
                {8'h2a,8'hxx,2'bx1} : dec_ma_data_saddr_op1 = 1'b1;  /* SUB,saddr,#byte */
                {8'h2b,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* SUB,A,saddr */
                {8'h3a,8'hxx,2'bx0} : dec_ma_data_saddr_op1 = 1'b1;  /* SUBC,saddr,#byte */
                {8'h3a,8'hxx,2'bx1} : dec_ma_data_saddr_op1 = 1'b1;  /* SUBC,saddr,#byte */
                {8'h3b,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* SUBC,A,saddr */
                {8'h5a,8'hxx,2'bx0} : dec_ma_data_saddr_op1 = 1'b1;  /* AND,saddr,#byte */
                {8'h5a,8'hxx,2'bx1} : dec_ma_data_saddr_op1 = 1'b1;  /* AND,saddr,#byte */
                {8'h5b,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* AND,A,saddr */
                {8'h6a,8'hxx,2'bx0} : dec_ma_data_saddr_op1 = 1'b1;  /* OR,saddr,#byte */
                {8'h6a,8'hxx,2'bx1} : dec_ma_data_saddr_op1 = 1'b1;  /* OR,saddr,#byte */
                {8'h6b,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* OR,A,saddr */
                {8'h7a,8'hxx,2'bx0} : dec_ma_data_saddr_op1 = 1'b1;  /* XOR,saddr,#byte */
                {8'h7a,8'hxx,2'bx1} : dec_ma_data_saddr_op1 = 1'b1;  /* XOR,saddr,#byte */
                {8'h7b,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* XOR,A,saddr */
                {8'h4a,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* CMP,saddr,#byte */
                {8'h4b,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* CMP,A,saddr */
                {8'hd4,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* CMP0,,saddr */
                {8'h06,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* ADDW,AX,saddrp */
                {8'h26,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* SUBW,AX,saddrp */
                {8'h46,8'hxx,2'bxx} : dec_ma_data_saddr_op1 = 1'b1;  /* CMPW,AX,saddrp */
                {8'ha4,8'hxx,2'bx0} : dec_ma_data_saddr_op1 = 1'b1;  /* INC,,saddr */
                {8'ha4,8'hxx,2'bx1} : dec_ma_data_saddr_op1 = 1'b1;  /* INC,,saddr */
                {8'hb4,8'hxx,2'bx0} : dec_ma_data_saddr_op1 = 1'b1;  /* DEC,,saddr */
                {8'hb4,8'hxx,2'bx1} : dec_ma_data_saddr_op1 = 1'b1;  /* DEC,,saddr */
                {8'ha6,8'hxx,2'bx0} : dec_ma_data_saddr_op1 = 1'b1;  /* INCW,,saddrp */
                {8'ha6,8'hxx,2'bx1} : dec_ma_data_saddr_op1 = 1'b1;  /* INCW,,saddrp */
                {8'hb6,8'hxx,2'bx0} : dec_ma_data_saddr_op1 = 1'b1;  /* DECW,,saddrp */
                {8'hb6,8'hxx,2'bx1} : dec_ma_data_saddr_op1 = 1'b1;  /* DECW,,saddrp */
                default : dec_ma_data_saddr_op1 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ma_data_saddr_op2;
    reg    dec_ma_data_saddr_op2;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_ma_data_saddr_op2 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hb8,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV,ES,saddr */
                {8'h61,8'ha8,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* XCH,A,saddr */
                {8'h61,8'ha8,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* XCH,A,saddr */
                {8'h71,8'h04,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,CY,saddr.0 */
                {8'h71,8'h14,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,CY,saddr.1 */
                {8'h71,8'h24,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,CY,saddr.2 */
                {8'h71,8'h34,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,CY,saddr.3 */
                {8'h71,8'h44,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,CY,saddr.4 */
                {8'h71,8'h54,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,CY,saddr.5 */
                {8'h71,8'h64,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,CY,saddr.6 */
                {8'h71,8'h74,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,CY,saddr.7 */
                {8'h71,8'h01,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,saddr.0,CY */
                {8'h71,8'h01,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,saddr.0,CY */
                {8'h71,8'h11,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,saddr.1,CY */
                {8'h71,8'h11,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,saddr.1,CY */
                {8'h71,8'h21,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,saddr.2,CY */
                {8'h71,8'h21,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,saddr.2,CY */
                {8'h71,8'h31,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,saddr.3,CY */
                {8'h71,8'h31,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,saddr.3,CY */
                {8'h71,8'h41,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,saddr.4,CY */
                {8'h71,8'h41,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,saddr.4,CY */
                {8'h71,8'h51,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,saddr.5,CY */
                {8'h71,8'h51,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,saddr.5,CY */
                {8'h71,8'h61,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,saddr.6,CY */
                {8'h71,8'h61,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,saddr.6,CY */
                {8'h71,8'h71,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,saddr.7,CY */
                {8'h71,8'h71,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* MOV1,saddr.7,CY */
                {8'h71,8'h05,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* AND1,CY,saddr.0 */
                {8'h71,8'h15,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* AND1,CY,saddr.1 */
                {8'h71,8'h25,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* AND1,CY,saddr.2 */
                {8'h71,8'h35,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* AND1,CY,saddr.3 */
                {8'h71,8'h45,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* AND1,CY,saddr.4 */
                {8'h71,8'h55,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* AND1,CY,saddr.5 */
                {8'h71,8'h65,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* AND1,CY,saddr.6 */
                {8'h71,8'h75,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* AND1,CY,saddr.7 */
                {8'h71,8'h06,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* OR1,CY,saddr.0 */
                {8'h71,8'h16,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* OR1,CY,saddr.1 */
                {8'h71,8'h26,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* OR1,CY,saddr.2 */
                {8'h71,8'h36,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* OR1,CY,saddr.3 */
                {8'h71,8'h46,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* OR1,CY,saddr.4 */
                {8'h71,8'h56,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* OR1,CY,saddr.5 */
                {8'h71,8'h66,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* OR1,CY,saddr.6 */
                {8'h71,8'h76,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* OR1,CY,saddr.7 */
                {8'h71,8'h07,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* XOR1,CY,saddr.0 */
                {8'h71,8'h17,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* XOR1,CY,saddr.1 */
                {8'h71,8'h27,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* XOR1,CY,saddr.2 */
                {8'h71,8'h37,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* XOR1,CY,saddr.3 */
                {8'h71,8'h47,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* XOR1,CY,saddr.4 */
                {8'h71,8'h57,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* XOR1,CY,saddr.5 */
                {8'h71,8'h67,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* XOR1,CY,saddr.6 */
                {8'h71,8'h77,2'bxx} : dec_ma_data_saddr_op2 = 1'b1;  /* XOR1,CY,saddr.7 */
                {8'h71,8'h02,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* SET1,,saddr.0 */
                {8'h71,8'h02,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* SET1,,saddr.0 */
                {8'h71,8'h12,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* SET1,,saddr.1 */
                {8'h71,8'h12,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* SET1,,saddr.1 */
                {8'h71,8'h22,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* SET1,,saddr.2 */
                {8'h71,8'h22,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* SET1,,saddr.2 */
                {8'h71,8'h32,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* SET1,,saddr.3 */
                {8'h71,8'h32,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* SET1,,saddr.3 */
                {8'h71,8'h42,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* SET1,,saddr.4 */
                {8'h71,8'h42,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* SET1,,saddr.4 */
                {8'h71,8'h52,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* SET1,,saddr.5 */
                {8'h71,8'h52,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* SET1,,saddr.5 */
                {8'h71,8'h62,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* SET1,,saddr.6 */
                {8'h71,8'h62,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* SET1,,saddr.6 */
                {8'h71,8'h72,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* SET1,,saddr.7 */
                {8'h71,8'h72,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* SET1,,saddr.7 */
                {8'h71,8'h03,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* CLR1,,saddr.0 */
                {8'h71,8'h03,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* CLR1,,saddr.0 */
                {8'h71,8'h13,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* CLR1,,saddr.1 */
                {8'h71,8'h13,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* CLR1,,saddr.1 */
                {8'h71,8'h23,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* CLR1,,saddr.2 */
                {8'h71,8'h23,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* CLR1,,saddr.2 */
                {8'h71,8'h33,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* CLR1,,saddr.3 */
                {8'h71,8'h33,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* CLR1,,saddr.3 */
                {8'h71,8'h43,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* CLR1,,saddr.4 */
                {8'h71,8'h43,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* CLR1,,saddr.4 */
                {8'h71,8'h53,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* CLR1,,saddr.5 */
                {8'h71,8'h53,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* CLR1,,saddr.5 */
                {8'h71,8'h63,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* CLR1,,saddr.6 */
                {8'h71,8'h63,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* CLR1,,saddr.6 */
                {8'h71,8'h73,2'bx0} : dec_ma_data_saddr_op2 = 1'b1;  /* CLR1,,saddr.7 */
                {8'h71,8'h73,2'bx1} : dec_ma_data_saddr_op2 = 1'b1;  /* CLR1,,saddr.7 */
                {8'h31,8'h02,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BT,saddr.0,$addr8 */
                {8'h31,8'h12,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BT,saddr.1,$addr8 */
                {8'h31,8'h22,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BT,saddr.2,$addr8 */
                {8'h31,8'h32,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BT,saddr.3,$addr8 */
                {8'h31,8'h42,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BT,saddr.4,$addr8 */
                {8'h31,8'h52,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BT,saddr.5,$addr8 */
                {8'h31,8'h62,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BT,saddr.6,$addr8 */
                {8'h31,8'h72,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BT,saddr.7,$addr8 */
                {8'h31,8'h04,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BF,saddr.0,$addr8 */
                {8'h31,8'h14,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BF,saddr.1,$addr8 */
                {8'h31,8'h24,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BF,saddr.2,$addr8 */
                {8'h31,8'h34,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BF,saddr.3,$addr8 */
                {8'h31,8'h44,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BF,saddr.4,$addr8 */
                {8'h31,8'h54,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BF,saddr.5,$addr8 */
                {8'h31,8'h64,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BF,saddr.6,$addr8 */
                {8'h31,8'h74,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BF,saddr.7,$addr8 */
                {8'h31,8'h00,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.0,$addr8 */
                {8'h31,8'h00,2'b01} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.0,$addr8 */
                {8'h31,8'h00,2'b10} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.0,$addr8 */
                {8'h31,8'h10,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.1,$addr8 */
                {8'h31,8'h10,2'b01} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.1,$addr8 */
                {8'h31,8'h10,2'b10} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.1,$addr8 */
                {8'h31,8'h20,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.2,$addr8 */
                {8'h31,8'h20,2'b01} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.2,$addr8 */
                {8'h31,8'h20,2'b10} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.2,$addr8 */
                {8'h31,8'h30,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.3,$addr8 */
                {8'h31,8'h30,2'b01} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.3,$addr8 */
                {8'h31,8'h30,2'b10} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.3,$addr8 */
                {8'h31,8'h40,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.4,$addr8 */
                {8'h31,8'h40,2'b01} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.4,$addr8 */
                {8'h31,8'h40,2'b10} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.4,$addr8 */
                {8'h31,8'h50,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.5,$addr8 */
                {8'h31,8'h50,2'b01} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.5,$addr8 */
                {8'h31,8'h50,2'b10} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.5,$addr8 */
                {8'h31,8'h60,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.6,$addr8 */
                {8'h31,8'h60,2'b01} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.6,$addr8 */
                {8'h31,8'h60,2'b10} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.6,$addr8 */
                {8'h31,8'h70,2'b00} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.7,$addr8 */
                {8'h31,8'h70,2'b01} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.7,$addr8 */
                {8'h31,8'h70,2'b10} : dec_ma_data_saddr_op2 = 1'b1;  /* BTCLR,saddr.7,$addr8 */
                default : dec_ma_data_saddr_op2 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ma_data_sfr_op1;
    reg    dec_ma_data_sfr_op1;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_ma_data_sfr_op1 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'hce,8'hxx,2'bxx} : dec_ma_data_sfr_op1 = 1'b1;  /* MOV,sfr,#byte */
                {8'h8e,8'hxx,2'bxx} : dec_ma_data_sfr_op1 = 1'b1;  /* MOV,A,sfr */
                {8'h9e,8'hxx,2'bxx} : dec_ma_data_sfr_op1 = 1'b1;  /* MOV,sfr,A */
                {8'hcb,8'hxx,2'bxx} : dec_ma_data_sfr_op1 = 1'b1;  /* MOVW,sfrp,#word */
                {8'hae,8'hxx,2'bxx} : dec_ma_data_sfr_op1 = 1'b1;  /* MOVW,AX,sfrp */
                {8'hbe,8'hxx,2'bxx} : dec_ma_data_sfr_op1 = 1'b1;  /* MOVW,sfrp,AX */
                default : dec_ma_data_sfr_op1 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ma_data_sfr_op2;
    reg    dec_ma_data_sfr_op2;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_ma_data_sfr_op2 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hab,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* XCH,A,sfr */
                {8'h61,8'hab,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* XCH,A,sfr */
                {8'h71,8'h0c,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,CY,sfr.0 */
                {8'h71,8'h1c,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,CY,sfr.1 */
                {8'h71,8'h2c,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,CY,sfr.2 */
                {8'h71,8'h3c,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,CY,sfr.3 */
                {8'h71,8'h4c,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,CY,sfr.4 */
                {8'h71,8'h5c,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,CY,sfr.5 */
                {8'h71,8'h6c,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,CY,sfr.6 */
                {8'h71,8'h7c,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,CY,sfr.7 */
                {8'h71,8'h09,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,sfr.0,CY */
                {8'h71,8'h09,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,sfr.0,CY */
                {8'h71,8'h19,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,sfr.1,CY */
                {8'h71,8'h19,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,sfr.1,CY */
                {8'h71,8'h29,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,sfr.2,CY */
                {8'h71,8'h29,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,sfr.2,CY */
                {8'h71,8'h39,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,sfr.3,CY */
                {8'h71,8'h39,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,sfr.3,CY */
                {8'h71,8'h49,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,sfr.4,CY */
                {8'h71,8'h49,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,sfr.4,CY */
                {8'h71,8'h59,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,sfr.5,CY */
                {8'h71,8'h59,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,sfr.5,CY */
                {8'h71,8'h69,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,sfr.6,CY */
                {8'h71,8'h69,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,sfr.6,CY */
                {8'h71,8'h79,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,sfr.7,CY */
                {8'h71,8'h79,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* MOV1,sfr.7,CY */
                {8'h71,8'h0d,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* AND1,CY,sfr.0 */
                {8'h71,8'h1d,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* AND1,CY,sfr.1 */
                {8'h71,8'h2d,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* AND1,CY,sfr.2 */
                {8'h71,8'h3d,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* AND1,CY,sfr.3 */
                {8'h71,8'h4d,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* AND1,CY,sfr.4 */
                {8'h71,8'h5d,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* AND1,CY,sfr.5 */
                {8'h71,8'h6d,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* AND1,CY,sfr.6 */
                {8'h71,8'h7d,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* AND1,CY,sfr.7 */
                {8'h71,8'h0e,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* OR1,CY,sfr.0 */
                {8'h71,8'h1e,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* OR1,CY,sfr.1 */
                {8'h71,8'h2e,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* OR1,CY,sfr.2 */
                {8'h71,8'h3e,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* OR1,CY,sfr.3 */
                {8'h71,8'h4e,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* OR1,CY,sfr.4 */
                {8'h71,8'h5e,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* OR1,CY,sfr.5 */
                {8'h71,8'h6e,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* OR1,CY,sfr.6 */
                {8'h71,8'h7e,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* OR1,CY,sfr.7 */
                {8'h71,8'h0f,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* XOR1,CY,sfr.0 */
                {8'h71,8'h1f,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* XOR1,CY,sfr.1 */
                {8'h71,8'h2f,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* XOR1,CY,sfr.2 */
                {8'h71,8'h3f,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* XOR1,CY,sfr.3 */
                {8'h71,8'h4f,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* XOR1,CY,sfr.4 */
                {8'h71,8'h5f,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* XOR1,CY,sfr.5 */
                {8'h71,8'h6f,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* XOR1,CY,sfr.6 */
                {8'h71,8'h7f,2'bxx} : dec_ma_data_sfr_op2 = 1'b1;  /* XOR1,CY,sfr.7 */
                {8'h71,8'h0a,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* SET1,,sfr.0 */
                {8'h71,8'h0a,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* SET1,,sfr.0 */
                {8'h71,8'h1a,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* SET1,,sfr.1 */
                {8'h71,8'h1a,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* SET1,,sfr.1 */
                {8'h71,8'h2a,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* SET1,,sfr.2 */
                {8'h71,8'h2a,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* SET1,,sfr.2 */
                {8'h71,8'h3a,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* SET1,,sfr.3 */
                {8'h71,8'h3a,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* SET1,,sfr.3 */
                {8'h71,8'h4a,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* SET1,,sfr.4 */
                {8'h71,8'h4a,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* SET1,,sfr.4 */
                {8'h71,8'h5a,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* SET1,,sfr.5 */
                {8'h71,8'h5a,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* SET1,,sfr.5 */
                {8'h71,8'h6a,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* SET1,,sfr.6 */
                {8'h71,8'h6a,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* SET1,,sfr.6 */
                {8'h71,8'h7a,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* SET1,,sfr.7 */
                {8'h71,8'h7a,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* SET1,,sfr.7 */
                {8'h71,8'h0b,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* CLR1,,sfr.0 */
                {8'h71,8'h0b,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* CLR1,,sfr.0 */
                {8'h71,8'h1b,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* CLR1,,sfr.1 */
                {8'h71,8'h1b,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* CLR1,,sfr.1 */
                {8'h71,8'h2b,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* CLR1,,sfr.2 */
                {8'h71,8'h2b,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* CLR1,,sfr.2 */
                {8'h71,8'h3b,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* CLR1,,sfr.3 */
                {8'h71,8'h3b,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* CLR1,,sfr.3 */
                {8'h71,8'h4b,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* CLR1,,sfr.4 */
                {8'h71,8'h4b,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* CLR1,,sfr.4 */
                {8'h71,8'h5b,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* CLR1,,sfr.5 */
                {8'h71,8'h5b,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* CLR1,,sfr.5 */
                {8'h71,8'h6b,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* CLR1,,sfr.6 */
                {8'h71,8'h6b,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* CLR1,,sfr.6 */
                {8'h71,8'h7b,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* CLR1,,sfr.7 */
                {8'h71,8'h7b,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* CLR1,,sfr.7 */
                {8'h31,8'h82,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BT,sfr.0,$addr8 */
                {8'h31,8'h92,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BT,sfr.1,$addr8 */
                {8'h31,8'ha2,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BT,sfr.2,$addr8 */
                {8'h31,8'hb2,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BT,sfr.3,$addr8 */
                {8'h31,8'hc2,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BT,sfr.4,$addr8 */
                {8'h31,8'hd2,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BT,sfr.5,$addr8 */
                {8'h31,8'he2,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BT,sfr.6,$addr8 */
                {8'h31,8'hf2,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BT,sfr.7,$addr8 */
                {8'h31,8'h84,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BF,sfr.0,$addr8 */
                {8'h31,8'h94,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BF,sfr.1,$addr8 */
                {8'h31,8'ha4,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BF,sfr.2,$addr8 */
                {8'h31,8'hb4,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BF,sfr.3,$addr8 */
                {8'h31,8'hc4,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BF,sfr.4,$addr8 */
                {8'h31,8'hd4,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BF,sfr.5,$addr8 */
                {8'h31,8'he4,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BF,sfr.6,$addr8 */
                {8'h31,8'hf4,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BF,sfr.7,$addr8 */
                {8'h31,8'h80,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.0,$addr8 */
                {8'h31,8'h80,2'b01} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.0,$addr8 */
                {8'h31,8'h80,2'b10} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.0,$addr8 */
                {8'h31,8'h90,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.1,$addr8 */
                {8'h31,8'h90,2'b01} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.1,$addr8 */
                {8'h31,8'h90,2'b10} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.1,$addr8 */
                {8'h31,8'ha0,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.2,$addr8 */
                {8'h31,8'ha0,2'b01} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.2,$addr8 */
                {8'h31,8'ha0,2'b10} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.2,$addr8 */
                {8'h31,8'hb0,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.3,$addr8 */
                {8'h31,8'hb0,2'b01} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.3,$addr8 */
                {8'h31,8'hb0,2'b10} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.3,$addr8 */
                {8'h31,8'hc0,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.4,$addr8 */
                {8'h31,8'hc0,2'b01} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.4,$addr8 */
                {8'h31,8'hc0,2'b10} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.4,$addr8 */
                {8'h31,8'hd0,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.5,$addr8 */
                {8'h31,8'hd0,2'b01} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.5,$addr8 */
                {8'h31,8'hd0,2'b10} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.5,$addr8 */
                {8'h31,8'he0,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.6,$addr8 */
                {8'h31,8'he0,2'b01} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.6,$addr8 */
                {8'h31,8'he0,2'b10} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.6,$addr8 */
                {8'h31,8'hf0,2'b00} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.7,$addr8 */
                {8'h31,8'hf0,2'b01} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.7,$addr8 */
                {8'h31,8'hf0,2'b10} : dec_ma_data_sfr_op2 = 1'b1;  /* BTCLR,sfr.7,$addr8 */
                {8'h61,8'hbb,2'bx0} : dec_ma_data_sfr_op2 = 1'b1;  /* XCH,A,sfr */
                {8'h61,8'hbb,2'bx1} : dec_ma_data_sfr_op2 = 1'b1;  /* XCH,A,sfr */
                default : dec_ma_data_sfr_op2 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ma_data_op12;
    reg    dec_ma_data_op12;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_ma_data_op12 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'hcf,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* MOV,!addr16,#byte */
                {8'h8f,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* MOV,A,!addr16 */
                {8'h9f,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* MOV,!addr16,A */
                {8'he9,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* MOV,B,!addr16 */
                {8'hf9,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* MOV,C,!addr16 */
                {8'hd9,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* MOV,X,!addr16 */
                {8'he5,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* ONEB,,!addr16 */
                {8'hf5,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* CLRB,,!addr16 */
                {8'haf,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* MOVW,AX,!addr16 */
                {8'hbf,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* MOVW,!addr16,AX */
                {8'hdb,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* MOVW,BC,!addr16 */
                {8'heb,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* MOVW,DE,!addr16 */
                {8'hfb,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* MOVW,HL,!addr16 */
                {8'h0f,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* ADD,A,!addr16 */
                {8'h1f,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* ADDC,A,!addr16 */
                {8'h2f,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* SUB,A,!addr16 */
                {8'h3f,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* SUBC,A,!addr16 */
                {8'h5f,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* AND,A,!addr16 */
                {8'h6f,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* OR,A,!addr16 */
                {8'h7f,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* XOR,A,!addr16 */
                {8'h40,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* CMP,!addr16,#byte */
                {8'h4f,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* CMP,A,!addr16 */
                {8'hd5,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* CMP0,,!addr16 */
                {8'h02,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* ADDW,AX,!addr16 */
                {8'h22,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* SUBW,AX,!addr16 */
                {8'h42,8'hxx,2'bxx} : dec_ma_data_op12 = 1'b1;  /* CMPW,AX,!addr16 */
                {8'ha0,8'hxx,2'bx0} : dec_ma_data_op12 = 1'b1;  /* INC,,!addr16 */
                {8'ha0,8'hxx,2'bx1} : dec_ma_data_op12 = 1'b1;  /* INC,,!addr16 */
                {8'hb0,8'hxx,2'bx0} : dec_ma_data_op12 = 1'b1;  /* DEC,,!addr16 */
                {8'hb0,8'hxx,2'bx1} : dec_ma_data_op12 = 1'b1;  /* DEC,,!addr16 */
                {8'ha2,8'hxx,2'bx0} : dec_ma_data_op12 = 1'b1;  /* INCW,,!addr16 */
                {8'ha2,8'hxx,2'bx1} : dec_ma_data_op12 = 1'b1;  /* INCW,,!addr16 */
                {8'hb2,8'hxx,2'bx0} : dec_ma_data_op12 = 1'b1;  /* DECW,,!addr16 */
                {8'hb2,8'hxx,2'bx1} : dec_ma_data_op12 = 1'b1;  /* DECW,,!addr16 */
                default : dec_ma_data_op12 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ma_data_op23;
    reg    dec_ma_data_op23;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_ma_data_op23 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'haa,2'bx0} : dec_ma_data_op23 = 1'b1;  /* XCH,A,!addr16 */
                {8'h61,8'haa,2'bx1} : dec_ma_data_op23 = 1'b1;  /* XCH,A,!addr16 */
                {8'h71,8'h00,2'bx0} : dec_ma_data_op23 = 1'b1;  /* SET1,,!addr16.0 */
                {8'h71,8'h00,2'bx1} : dec_ma_data_op23 = 1'b1;  /* SET1,,!addr16.0 */
                {8'h71,8'h10,2'bx0} : dec_ma_data_op23 = 1'b1;  /* SET1,,!addr16.1 */
                {8'h71,8'h10,2'bx1} : dec_ma_data_op23 = 1'b1;  /* SET1,,!addr16.1 */
                {8'h71,8'h20,2'bx0} : dec_ma_data_op23 = 1'b1;  /* SET1,,!addr16.2 */
                {8'h71,8'h20,2'bx1} : dec_ma_data_op23 = 1'b1;  /* SET1,,!addr16.2 */
                {8'h71,8'h30,2'bx0} : dec_ma_data_op23 = 1'b1;  /* SET1,,!addr16.3 */
                {8'h71,8'h30,2'bx1} : dec_ma_data_op23 = 1'b1;  /* SET1,,!addr16.3 */
                {8'h71,8'h40,2'bx0} : dec_ma_data_op23 = 1'b1;  /* SET1,,!addr16.4 */
                {8'h71,8'h40,2'bx1} : dec_ma_data_op23 = 1'b1;  /* SET1,,!addr16.4 */
                {8'h71,8'h50,2'bx0} : dec_ma_data_op23 = 1'b1;  /* SET1,,!addr16.5 */
                {8'h71,8'h50,2'bx1} : dec_ma_data_op23 = 1'b1;  /* SET1,,!addr16.5 */
                {8'h71,8'h60,2'bx0} : dec_ma_data_op23 = 1'b1;  /* SET1,,!addr16.6 */
                {8'h71,8'h60,2'bx1} : dec_ma_data_op23 = 1'b1;  /* SET1,,!addr16.6 */
                {8'h71,8'h70,2'bx0} : dec_ma_data_op23 = 1'b1;  /* SET1,,!addr16.7 */
                {8'h71,8'h70,2'bx1} : dec_ma_data_op23 = 1'b1;  /* SET1,,!addr16.7 */
                {8'h71,8'h08,2'bx0} : dec_ma_data_op23 = 1'b1;  /* CLR1,,!addr16.0 */
                {8'h71,8'h08,2'bx1} : dec_ma_data_op23 = 1'b1;  /* CLR1,,!addr16.0 */
                {8'h71,8'h18,2'bx0} : dec_ma_data_op23 = 1'b1;  /* CLR1,,!addr16.1 */
                {8'h71,8'h18,2'bx1} : dec_ma_data_op23 = 1'b1;  /* CLR1,,!addr16.1 */
                {8'h71,8'h28,2'bx0} : dec_ma_data_op23 = 1'b1;  /* CLR1,,!addr16.2 */
                {8'h71,8'h28,2'bx1} : dec_ma_data_op23 = 1'b1;  /* CLR1,,!addr16.2 */
                {8'h71,8'h38,2'bx0} : dec_ma_data_op23 = 1'b1;  /* CLR1,,!addr16.3 */
                {8'h71,8'h38,2'bx1} : dec_ma_data_op23 = 1'b1;  /* CLR1,,!addr16.3 */
                {8'h71,8'h48,2'bx0} : dec_ma_data_op23 = 1'b1;  /* CLR1,,!addr16.4 */
                {8'h71,8'h48,2'bx1} : dec_ma_data_op23 = 1'b1;  /* CLR1,,!addr16.4 */
                {8'h71,8'h58,2'bx0} : dec_ma_data_op23 = 1'b1;  /* CLR1,,!addr16.5 */
                {8'h71,8'h58,2'bx1} : dec_ma_data_op23 = 1'b1;  /* CLR1,,!addr16.5 */
                {8'h71,8'h68,2'bx0} : dec_ma_data_op23 = 1'b1;  /* CLR1,,!addr16.6 */
                {8'h71,8'h68,2'bx1} : dec_ma_data_op23 = 1'b1;  /* CLR1,,!addr16.6 */
                {8'h71,8'h78,2'bx0} : dec_ma_data_op23 = 1'b1;  /* CLR1,,!addr16.7 */
                {8'h71,8'h78,2'bx1} : dec_ma_data_op23 = 1'b1;  /* CLR1,,!addr16.7 */
                {8'h61,8'hba,2'bx0} : dec_ma_data_op23 = 1'b1;  /* XCH,A,!addr16 */
                {8'h61,8'hba,2'bx1} : dec_ma_data_op23 = 1'b1;  /* XCH,A,!addr16 */
                default : dec_ma_data_op23 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ma_data_HL;
    reg    dec_ma_data_HL;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_ma_data_HL = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h8b,8'hxx,2'bxx} : dec_ma_data_HL = 1'b1;  /* MOV,A,[HL] */
                {8'h9b,8'hxx,2'bxx} : dec_ma_data_HL = 1'b1;  /* MOV,[HL],A */
                {8'h61,8'hac,2'bx0} : dec_ma_data_HL = 1'b1;  /* XCH,A,[HL] */
                {8'h61,8'hac,2'bx1} : dec_ma_data_HL = 1'b1;  /* XCH,A,[HL] */
                {8'hab,8'hxx,2'bxx} : dec_ma_data_HL = 1'b1;  /* MOVW,AX,[HL] */
                {8'hbb,8'hxx,2'bxx} : dec_ma_data_HL = 1'b1;  /* MOVW,[HL],AX */
                {8'h0d,8'hxx,2'bxx} : dec_ma_data_HL = 1'b1;  /* ADD,A,[HL] */
                {8'h1d,8'hxx,2'bxx} : dec_ma_data_HL = 1'b1;  /* ADDC,A,[HL] */
                {8'h2d,8'hxx,2'bxx} : dec_ma_data_HL = 1'b1;  /* SUB,A,[HL] */
                {8'h3d,8'hxx,2'bxx} : dec_ma_data_HL = 1'b1;  /* SUBC,A,[HL] */
                {8'h5d,8'hxx,2'bxx} : dec_ma_data_HL = 1'b1;  /* AND,A,[HL] */
                {8'h6d,8'hxx,2'bxx} : dec_ma_data_HL = 1'b1;  /* OR,A,[HL] */
                {8'h7d,8'hxx,2'bxx} : dec_ma_data_HL = 1'b1;  /* XOR,A,[HL] */
                {8'h4d,8'hxx,2'bxx} : dec_ma_data_HL = 1'b1;  /* CMP,A,[HL] */
                {8'h71,8'h84,2'bxx} : dec_ma_data_HL = 1'b1;  /* MOV1,CY,[HL].0 */
                {8'h71,8'h94,2'bxx} : dec_ma_data_HL = 1'b1;  /* MOV1,CY,[HL].1 */
                {8'h71,8'ha4,2'bxx} : dec_ma_data_HL = 1'b1;  /* MOV1,CY,[HL].2 */
                {8'h71,8'hb4,2'bxx} : dec_ma_data_HL = 1'b1;  /* MOV1,CY,[HL].3 */
                {8'h71,8'hc4,2'bxx} : dec_ma_data_HL = 1'b1;  /* MOV1,CY,[HL].4 */
                {8'h71,8'hd4,2'bxx} : dec_ma_data_HL = 1'b1;  /* MOV1,CY,[HL].5 */
                {8'h71,8'he4,2'bxx} : dec_ma_data_HL = 1'b1;  /* MOV1,CY,[HL].6 */
                {8'h71,8'hf4,2'bxx} : dec_ma_data_HL = 1'b1;  /* MOV1,CY,[HL].7 */
                {8'h71,8'h81,2'bx0} : dec_ma_data_HL = 1'b1;  /* MOV1,[HL].0,CY */
                {8'h71,8'h81,2'bx1} : dec_ma_data_HL = 1'b1;  /* MOV1,[HL].0,CY */
                {8'h71,8'h91,2'bx0} : dec_ma_data_HL = 1'b1;  /* MOV1,[HL].1,CY */
                {8'h71,8'h91,2'bx1} : dec_ma_data_HL = 1'b1;  /* MOV1,[HL].1,CY */
                {8'h71,8'ha1,2'bx0} : dec_ma_data_HL = 1'b1;  /* MOV1,[HL].2,CY */
                {8'h71,8'ha1,2'bx1} : dec_ma_data_HL = 1'b1;  /* MOV1,[HL].2,CY */
                {8'h71,8'hb1,2'bx0} : dec_ma_data_HL = 1'b1;  /* MOV1,[HL].3,CY */
                {8'h71,8'hb1,2'bx1} : dec_ma_data_HL = 1'b1;  /* MOV1,[HL].3,CY */
                {8'h71,8'hc1,2'bx0} : dec_ma_data_HL = 1'b1;  /* MOV1,[HL].4,CY */
                {8'h71,8'hc1,2'bx1} : dec_ma_data_HL = 1'b1;  /* MOV1,[HL].4,CY */
                {8'h71,8'hd1,2'bx0} : dec_ma_data_HL = 1'b1;  /* MOV1,[HL].5,CY */
                {8'h71,8'hd1,2'bx1} : dec_ma_data_HL = 1'b1;  /* MOV1,[HL].5,CY */
                {8'h71,8'he1,2'bx0} : dec_ma_data_HL = 1'b1;  /* MOV1,[HL].6,CY */
                {8'h71,8'he1,2'bx1} : dec_ma_data_HL = 1'b1;  /* MOV1,[HL].6,CY */
                {8'h71,8'hf1,2'bx0} : dec_ma_data_HL = 1'b1;  /* MOV1,[HL].7,CY */
                {8'h71,8'hf1,2'bx1} : dec_ma_data_HL = 1'b1;  /* MOV1,[HL].7,CY */
                {8'h71,8'h85,2'bxx} : dec_ma_data_HL = 1'b1;  /* AND1,CY,[HL].0 */
                {8'h71,8'h95,2'bxx} : dec_ma_data_HL = 1'b1;  /* AND1,CY,[HL].1 */
                {8'h71,8'ha5,2'bxx} : dec_ma_data_HL = 1'b1;  /* AND1,CY,[HL].2 */
                {8'h71,8'hb5,2'bxx} : dec_ma_data_HL = 1'b1;  /* AND1,CY,[HL].3 */
                {8'h71,8'hc5,2'bxx} : dec_ma_data_HL = 1'b1;  /* AND1,CY,[HL].4 */
                {8'h71,8'hd5,2'bxx} : dec_ma_data_HL = 1'b1;  /* AND1,CY,[HL].5 */
                {8'h71,8'he5,2'bxx} : dec_ma_data_HL = 1'b1;  /* AND1,CY,[HL].6 */
                {8'h71,8'hf5,2'bxx} : dec_ma_data_HL = 1'b1;  /* AND1,CY,[HL].7 */
                {8'h71,8'h86,2'bxx} : dec_ma_data_HL = 1'b1;  /* OR1,CY,[HL].0 */
                {8'h71,8'h96,2'bxx} : dec_ma_data_HL = 1'b1;  /* OR1,CY,[HL].1 */
                {8'h71,8'ha6,2'bxx} : dec_ma_data_HL = 1'b1;  /* OR1,CY,[HL].2 */
                {8'h71,8'hb6,2'bxx} : dec_ma_data_HL = 1'b1;  /* OR1,CY,[HL].3 */
                {8'h71,8'hc6,2'bxx} : dec_ma_data_HL = 1'b1;  /* OR1,CY,[HL].4 */
                {8'h71,8'hd6,2'bxx} : dec_ma_data_HL = 1'b1;  /* OR1,CY,[HL].5 */
                {8'h71,8'he6,2'bxx} : dec_ma_data_HL = 1'b1;  /* OR1,CY,[HL].6 */
                {8'h71,8'hf6,2'bxx} : dec_ma_data_HL = 1'b1;  /* OR1,CY,[HL].7 */
                {8'h71,8'h87,2'bxx} : dec_ma_data_HL = 1'b1;  /* XOR1,CY,[HL].0 */
                {8'h71,8'h97,2'bxx} : dec_ma_data_HL = 1'b1;  /* XOR1,CY,[HL].1 */
                {8'h71,8'ha7,2'bxx} : dec_ma_data_HL = 1'b1;  /* XOR1,CY,[HL].2 */
                {8'h71,8'hb7,2'bxx} : dec_ma_data_HL = 1'b1;  /* XOR1,CY,[HL].3 */
                {8'h71,8'hc7,2'bxx} : dec_ma_data_HL = 1'b1;  /* XOR1,CY,[HL].4 */
                {8'h71,8'hd7,2'bxx} : dec_ma_data_HL = 1'b1;  /* XOR1,CY,[HL].5 */
                {8'h71,8'he7,2'bxx} : dec_ma_data_HL = 1'b1;  /* XOR1,CY,[HL].6 */
                {8'h71,8'hf7,2'bxx} : dec_ma_data_HL = 1'b1;  /* XOR1,CY,[HL].7 */
                {8'h71,8'h82,2'bx0} : dec_ma_data_HL = 1'b1;  /* SET1,,[HL].0 */
                {8'h71,8'h82,2'bx1} : dec_ma_data_HL = 1'b1;  /* SET1,,[HL].0 */
                {8'h71,8'h92,2'bx0} : dec_ma_data_HL = 1'b1;  /* SET1,,[HL].1 */
                {8'h71,8'h92,2'bx1} : dec_ma_data_HL = 1'b1;  /* SET1,,[HL].1 */
                {8'h71,8'ha2,2'bx0} : dec_ma_data_HL = 1'b1;  /* SET1,,[HL].2 */
                {8'h71,8'ha2,2'bx1} : dec_ma_data_HL = 1'b1;  /* SET1,,[HL].2 */
                {8'h71,8'hb2,2'bx0} : dec_ma_data_HL = 1'b1;  /* SET1,,[HL].3 */
                {8'h71,8'hb2,2'bx1} : dec_ma_data_HL = 1'b1;  /* SET1,,[HL].3 */
                {8'h71,8'hc2,2'bx0} : dec_ma_data_HL = 1'b1;  /* SET1,,[HL].4 */
                {8'h71,8'hc2,2'bx1} : dec_ma_data_HL = 1'b1;  /* SET1,,[HL].4 */
                {8'h71,8'hd2,2'bx0} : dec_ma_data_HL = 1'b1;  /* SET1,,[HL].5 */
                {8'h71,8'hd2,2'bx1} : dec_ma_data_HL = 1'b1;  /* SET1,,[HL].5 */
                {8'h71,8'he2,2'bx0} : dec_ma_data_HL = 1'b1;  /* SET1,,[HL].6 */
                {8'h71,8'he2,2'bx1} : dec_ma_data_HL = 1'b1;  /* SET1,,[HL].6 */
                {8'h71,8'hf2,2'bx0} : dec_ma_data_HL = 1'b1;  /* SET1,,[HL].7 */
                {8'h71,8'hf2,2'bx1} : dec_ma_data_HL = 1'b1;  /* SET1,,[HL].7 */
                {8'h71,8'h83,2'bx0} : dec_ma_data_HL = 1'b1;  /* CLR1,,[HL].0 */
                {8'h71,8'h83,2'bx1} : dec_ma_data_HL = 1'b1;  /* CLR1,,[HL].0 */
                {8'h71,8'h93,2'bx0} : dec_ma_data_HL = 1'b1;  /* CLR1,,[HL].1 */
                {8'h71,8'h93,2'bx1} : dec_ma_data_HL = 1'b1;  /* CLR1,,[HL].1 */
                {8'h71,8'ha3,2'bx0} : dec_ma_data_HL = 1'b1;  /* CLR1,,[HL].2 */
                {8'h71,8'ha3,2'bx1} : dec_ma_data_HL = 1'b1;  /* CLR1,,[HL].2 */
                {8'h71,8'hb3,2'bx0} : dec_ma_data_HL = 1'b1;  /* CLR1,,[HL].3 */
                {8'h71,8'hb3,2'bx1} : dec_ma_data_HL = 1'b1;  /* CLR1,,[HL].3 */
                {8'h71,8'hc3,2'bx0} : dec_ma_data_HL = 1'b1;  /* CLR1,,[HL].4 */
                {8'h71,8'hc3,2'bx1} : dec_ma_data_HL = 1'b1;  /* CLR1,,[HL].4 */
                {8'h71,8'hd3,2'bx0} : dec_ma_data_HL = 1'b1;  /* CLR1,,[HL].5 */
                {8'h71,8'hd3,2'bx1} : dec_ma_data_HL = 1'b1;  /* CLR1,,[HL].5 */
                {8'h71,8'he3,2'bx0} : dec_ma_data_HL = 1'b1;  /* CLR1,,[HL].6 */
                {8'h71,8'he3,2'bx1} : dec_ma_data_HL = 1'b1;  /* CLR1,,[HL].6 */
                {8'h71,8'hf3,2'bx0} : dec_ma_data_HL = 1'b1;  /* CLR1,,[HL].7 */
                {8'h71,8'hf3,2'bx1} : dec_ma_data_HL = 1'b1;  /* CLR1,,[HL].7 */
                {8'h31,8'h83,2'b00} : dec_ma_data_HL = 1'b1;  /* BT,[HL].0,$addr8 */
                {8'h31,8'h93,2'b00} : dec_ma_data_HL = 1'b1;  /* BT,[HL].1,$addr8 */
                {8'h31,8'ha3,2'b00} : dec_ma_data_HL = 1'b1;  /* BT,[HL].2,$addr8 */
                {8'h31,8'hb3,2'b00} : dec_ma_data_HL = 1'b1;  /* BT,[HL].3,$addr8 */
                {8'h31,8'hc3,2'b00} : dec_ma_data_HL = 1'b1;  /* BT,[HL].4,$addr8 */
                {8'h31,8'hd3,2'b00} : dec_ma_data_HL = 1'b1;  /* BT,[HL].5,$addr8 */
                {8'h31,8'he3,2'b00} : dec_ma_data_HL = 1'b1;  /* BT,[HL].6,$addr8 */
                {8'h31,8'hf3,2'b00} : dec_ma_data_HL = 1'b1;  /* BT,[HL].7,$addr8 */
                {8'h31,8'h85,2'b00} : dec_ma_data_HL = 1'b1;  /* BF,[HL].0,$addr8 */
                {8'h31,8'h95,2'b00} : dec_ma_data_HL = 1'b1;  /* BF,[HL].1,$addr8 */
                {8'h31,8'ha5,2'b00} : dec_ma_data_HL = 1'b1;  /* BF,[HL].2,$addr8 */
                {8'h31,8'hb5,2'b00} : dec_ma_data_HL = 1'b1;  /* BF,[HL].3,$addr8 */
                {8'h31,8'hc5,2'b00} : dec_ma_data_HL = 1'b1;  /* BF,[HL].4,$addr8 */
                {8'h31,8'hd5,2'b00} : dec_ma_data_HL = 1'b1;  /* BF,[HL].5,$addr8 */
                {8'h31,8'he5,2'b00} : dec_ma_data_HL = 1'b1;  /* BF,[HL].6,$addr8 */
                {8'h31,8'hf5,2'b00} : dec_ma_data_HL = 1'b1;  /* BF,[HL].7,$addr8 */
                {8'h31,8'h81,2'b00} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].0,$addr8 */
                {8'h31,8'h81,2'b01} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].0,$addr8 */
                {8'h31,8'h81,2'b10} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].0,$addr8 */
                {8'h31,8'h91,2'b00} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].1,$addr8 */
                {8'h31,8'h91,2'b01} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].1,$addr8 */
                {8'h31,8'h91,2'b10} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].1,$addr8 */
                {8'h31,8'ha1,2'b00} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].2,$addr8 */
                {8'h31,8'ha1,2'b01} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].2,$addr8 */
                {8'h31,8'ha1,2'b10} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].2,$addr8 */
                {8'h31,8'hb1,2'b00} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].3,$addr8 */
                {8'h31,8'hb1,2'b01} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].3,$addr8 */
                {8'h31,8'hb1,2'b10} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].3,$addr8 */
                {8'h31,8'hc1,2'b00} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].4,$addr8 */
                {8'h31,8'hc1,2'b01} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].4,$addr8 */
                {8'h31,8'hc1,2'b10} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].4,$addr8 */
                {8'h31,8'hd1,2'b00} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].5,$addr8 */
                {8'h31,8'hd1,2'b01} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].5,$addr8 */
                {8'h31,8'hd1,2'b10} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].5,$addr8 */
                {8'h31,8'he1,2'b00} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].6,$addr8 */
                {8'h31,8'he1,2'b01} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].6,$addr8 */
                {8'h31,8'he1,2'b10} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].6,$addr8 */
                {8'h31,8'hf1,2'b00} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].7,$addr8 */
                {8'h31,8'hf1,2'b01} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].7,$addr8 */
                {8'h31,8'hf1,2'b10} : dec_ma_data_HL = 1'b1;  /* BTCLR,[HL].7,$addr8 */
                {8'h61,8'hbc,2'bx0} : dec_ma_data_HL = 1'b1;  /* XCH,A,[HL] */
                {8'h61,8'hbc,2'bx1} : dec_ma_data_HL = 1'b1;  /* XCH,A,[HL] */
                default : dec_ma_data_HL = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ma_data_HLop1;
    reg    dec_ma_data_HLop1;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_ma_data_HLop1 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'hcc,8'hxx,2'bxx} : dec_ma_data_HLop1 = 1'b1;  /* MOV,[HL+byte],#byte */
                {8'h8c,8'hxx,2'bxx} : dec_ma_data_HLop1 = 1'b1;  /* MOV,A,[HL+byte] */
                {8'h9c,8'hxx,2'bxx} : dec_ma_data_HLop1 = 1'b1;  /* MOV,[HL+byte],A */
                {8'hac,8'hxx,2'bxx} : dec_ma_data_HLop1 = 1'b1;  /* MOVW,AX,[HL+byte] */
                {8'hbc,8'hxx,2'bxx} : dec_ma_data_HLop1 = 1'b1;  /* MOVW,[HL+byte],AX */
                {8'h0e,8'hxx,2'bxx} : dec_ma_data_HLop1 = 1'b1;  /* ADD,A,[HL+byte] */
                {8'h1e,8'hxx,2'bxx} : dec_ma_data_HLop1 = 1'b1;  /* ADDC,A,[HL+byte] */
                {8'h2e,8'hxx,2'bxx} : dec_ma_data_HLop1 = 1'b1;  /* SUB,A,[HL+byte] */
                {8'h3e,8'hxx,2'bxx} : dec_ma_data_HLop1 = 1'b1;  /* SUBC,A,[HL+byte] */
                {8'h5e,8'hxx,2'bxx} : dec_ma_data_HLop1 = 1'b1;  /* AND,A,[HL+byte] */
                {8'h6e,8'hxx,2'bxx} : dec_ma_data_HLop1 = 1'b1;  /* OR,A,[HL+byte] */
                {8'h7e,8'hxx,2'bxx} : dec_ma_data_HLop1 = 1'b1;  /* XOR,A,[HL+byte] */
                {8'h4e,8'hxx,2'bxx} : dec_ma_data_HLop1 = 1'b1;  /* CMP,A,[HL+byte] */
                default : dec_ma_data_HLop1 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ma_data_HLop2;
    reg    dec_ma_data_HLop2;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_ma_data_HLop2 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hce,2'bxx} : dec_ma_data_HLop2 = 1'b1;  /* MOVS,[HL+byte],X */
                {8'h61,8'had,2'bx0} : dec_ma_data_HLop2 = 1'b1;  /* XCH,A,[HL+byte] */
                {8'h61,8'had,2'bx1} : dec_ma_data_HLop2 = 1'b1;  /* XCH,A,[HL+byte] */
                {8'h61,8'hde,2'bxx} : dec_ma_data_HLop2 = 1'b1;  /* CMPS,X,[HL+byte] */
                {8'h61,8'h09,2'bxx} : dec_ma_data_HLop2 = 1'b1;  /* ADDW,AX,[HL+byte] */
                {8'h61,8'h29,2'bxx} : dec_ma_data_HLop2 = 1'b1;  /* SUBW,AX,[HL+byte] */
                {8'h61,8'h49,2'bxx} : dec_ma_data_HLop2 = 1'b1;  /* CMPW,AX,[HL+byte] */
                {8'h61,8'h59,2'bx0} : dec_ma_data_HLop2 = 1'b1;  /* INC,,[HL+byte] */
                {8'h61,8'h59,2'bx1} : dec_ma_data_HLop2 = 1'b1;  /* INC,,[HL+byte] */
                {8'h61,8'h69,2'bx0} : dec_ma_data_HLop2 = 1'b1;  /* DEC,,[HL+byte] */
                {8'h61,8'h69,2'bx1} : dec_ma_data_HLop2 = 1'b1;  /* DEC,,[HL+byte] */
                {8'h61,8'h79,2'bx0} : dec_ma_data_HLop2 = 1'b1;  /* INCW,,[HL+byte] */
                {8'h61,8'h79,2'bx1} : dec_ma_data_HLop2 = 1'b1;  /* INCW,,[HL+byte] */
                {8'h61,8'h89,2'bx0} : dec_ma_data_HLop2 = 1'b1;  /* DECW,,[HL+byte] */
                {8'h61,8'h89,2'bx1} : dec_ma_data_HLop2 = 1'b1;  /* DECW,,[HL+byte] */
                {8'h61,8'hbd,2'bx0} : dec_ma_data_HLop2 = 1'b1;  /* XCH,A,[HL+byte] */
                {8'h61,8'hbd,2'bx1} : dec_ma_data_HLop2 = 1'b1;  /* XCH,A,[HL+byte] */
                default : dec_ma_data_HLop2 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ma_data_HLB;
    reg    dec_ma_data_HLB;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_ma_data_HLB = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hc9,2'bxx} : dec_ma_data_HLB = 1'b1;  /* MOV,A,[HL+B] */
                {8'h61,8'hd9,2'bxx} : dec_ma_data_HLB = 1'b1;  /* MOV,[HL+B],A */
                {8'h61,8'hb9,2'bx0} : dec_ma_data_HLB = 1'b1;  /* XCH,A,[HL+B] */
                {8'h61,8'hb9,2'bx1} : dec_ma_data_HLB = 1'b1;  /* XCH,A,[HL+B] */
                {8'h61,8'h80,2'bxx} : dec_ma_data_HLB = 1'b1;  /* ADD,A,[HL+B] */
                {8'h61,8'h90,2'bxx} : dec_ma_data_HLB = 1'b1;  /* ADDC,A,[HL+B] */
                {8'h61,8'ha0,2'bxx} : dec_ma_data_HLB = 1'b1;  /* SUB,A,[HL+B] */
                {8'h61,8'hb0,2'bxx} : dec_ma_data_HLB = 1'b1;  /* SUBC,A,[HL+B] */
                {8'h61,8'hd0,2'bxx} : dec_ma_data_HLB = 1'b1;  /* AND,A,[HL+B] */
                {8'h61,8'he0,2'bxx} : dec_ma_data_HLB = 1'b1;  /* OR,A,[HL+B] */
                {8'h61,8'hf0,2'bxx} : dec_ma_data_HLB = 1'b1;  /* XOR,A,[HL+B] */
                {8'h61,8'hc0,2'bxx} : dec_ma_data_HLB = 1'b1;  /* CMP,A,[HL+B] */
                {8'h61,8'hd1,2'bxx} : dec_ma_data_HLB = 1'b1;  /* AND,A,[HL+B] */
                {8'h61,8'he1,2'bxx} : dec_ma_data_HLB = 1'b1;  /* OR,A,[HL+B] */
                {8'h61,8'hf1,2'bxx} : dec_ma_data_HLB = 1'b1;  /* XOR,A,[HL+B] */
                default : dec_ma_data_HLB = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ma_data_HLC;
    reg    dec_ma_data_HLC;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_ma_data_HLC = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'he9,2'bxx} : dec_ma_data_HLC = 1'b1;  /* MOV,A,[HL+C] */
                {8'h61,8'hf9,2'bxx} : dec_ma_data_HLC = 1'b1;  /* MOV,[HL+C],A */
                {8'h61,8'ha9,2'bx0} : dec_ma_data_HLC = 1'b1;  /* XCH,A,[HL+C] */
                {8'h61,8'ha9,2'bx1} : dec_ma_data_HLC = 1'b1;  /* XCH,A,[HL+C] */
                {8'h61,8'h82,2'bxx} : dec_ma_data_HLC = 1'b1;  /* ADD,A,[HL+C] */
                {8'h61,8'h92,2'bxx} : dec_ma_data_HLC = 1'b1;  /* ADDC,A,[HL+C] */
                {8'h61,8'ha2,2'bxx} : dec_ma_data_HLC = 1'b1;  /* SUB,A,[HL+C] */
                {8'h61,8'hb2,2'bxx} : dec_ma_data_HLC = 1'b1;  /* SUBC,A,[HL+C] */
                {8'h61,8'hd2,2'bxx} : dec_ma_data_HLC = 1'b1;  /* AND,A,[HL+C] */
                {8'h61,8'he2,2'bxx} : dec_ma_data_HLC = 1'b1;  /* OR,A,[HL+C] */
                {8'h61,8'hf2,2'bxx} : dec_ma_data_HLC = 1'b1;  /* XOR,A,[HL+C] */
                {8'h61,8'hc2,2'bxx} : dec_ma_data_HLC = 1'b1;  /* CMP,A,[HL+C] */
                {8'h61,8'h83,2'bxx} : dec_ma_data_HLC = 1'b1;  /* ADD,A,[HL+C] */
                {8'h61,8'h93,2'bxx} : dec_ma_data_HLC = 1'b1;  /* ADDC,A,[HL+C] */
                {8'h61,8'ha3,2'bxx} : dec_ma_data_HLC = 1'b1;  /* SUB,A,[HL+C] */
                {8'h61,8'hb3,2'bxx} : dec_ma_data_HLC = 1'b1;  /* SUBC,A,[HL+C] */
                default : dec_ma_data_HLC = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ma_data_DE;
    reg    dec_ma_data_DE;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_ma_data_DE = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h89,8'hxx,2'bxx} : dec_ma_data_DE = 1'b1;  /* MOV,A,[DE] */
                {8'h99,8'hxx,2'bxx} : dec_ma_data_DE = 1'b1;  /* MOV,[DE],A */
                {8'h61,8'hae,2'bx0} : dec_ma_data_DE = 1'b1;  /* XCH,A,[DE] */
                {8'h61,8'hae,2'bx1} : dec_ma_data_DE = 1'b1;  /* XCH,A,[DE] */
                {8'ha9,8'hxx,2'bxx} : dec_ma_data_DE = 1'b1;  /* MOVW,AX,[DE] */
                {8'hb9,8'hxx,2'bxx} : dec_ma_data_DE = 1'b1;  /* MOVW,[DE],AX */
                {8'h61,8'hbe,2'bx0} : dec_ma_data_DE = 1'b1;  /* XCH,A,[DE] */
                {8'h61,8'hbe,2'bx1} : dec_ma_data_DE = 1'b1;  /* XCH,A,[DE] */
                default : dec_ma_data_DE = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ma_data_DEop1;
    reg    dec_ma_data_DEop1;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_ma_data_DEop1 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'hca,8'hxx,2'bxx} : dec_ma_data_DEop1 = 1'b1;  /* MOV,[DE+byte],#byte */
                {8'h8a,8'hxx,2'bxx} : dec_ma_data_DEop1 = 1'b1;  /* MOV,A,[DE+byte] */
                {8'h9a,8'hxx,2'bxx} : dec_ma_data_DEop1 = 1'b1;  /* MOV,[DE+byte],A */
                {8'haa,8'hxx,2'bxx} : dec_ma_data_DEop1 = 1'b1;  /* MOVW,AX,[DE+byte] */
                {8'hba,8'hxx,2'bxx} : dec_ma_data_DEop1 = 1'b1;  /* MOVW,[DE+byte],AX */
                default : dec_ma_data_DEop1 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ma_data_DEop2;
    reg    dec_ma_data_DEop2;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_ma_data_DEop2 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'haf,2'bx0} : dec_ma_data_DEop2 = 1'b1;  /* XCH,A,[DE+byte] */
                {8'h61,8'haf,2'bx1} : dec_ma_data_DEop2 = 1'b1;  /* XCH,A,[DE+byte] */
                {8'h61,8'hbf,2'bx0} : dec_ma_data_DEop2 = 1'b1;  /* XCH,A,[DE+byte] */
                {8'h61,8'hbf,2'bx1} : dec_ma_data_DEop2 = 1'b1;  /* XCH,A,[DE+byte] */
                default : dec_ma_data_DEop2 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ma_data_SPop1;
    reg    dec_ma_data_SPop1;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_ma_data_SPop1 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'hc8,8'hxx,2'bxx} : dec_ma_data_SPop1 = 1'b1;  /* MOV,[SP+byte],#byte */
                {8'h88,8'hxx,2'bxx} : dec_ma_data_SPop1 = 1'b1;  /* MOV,A,[SP+byte] */
                {8'h98,8'hxx,2'bxx} : dec_ma_data_SPop1 = 1'b1;  /* MOV,[SP+byte],A */
                {8'ha8,8'hxx,2'bxx} : dec_ma_data_SPop1 = 1'b1;  /* MOVW,AX,[SP+byte] */
                {8'hb8,8'hxx,2'bxx} : dec_ma_data_SPop1 = 1'b1;  /* MOVW,[SP+byte],AX */
                default : dec_ma_data_SPop1 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ma_data_BCop12;
    reg    dec_ma_data_BCop12;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_ma_data_BCop12 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h39,8'hxx,2'bxx} : dec_ma_data_BCop12 = 1'b1;  /* MOV,word[BC],#byte */
                {8'h49,8'hxx,2'bxx} : dec_ma_data_BCop12 = 1'b1;  /* MOV,A,word[BC] */
                {8'h48,8'hxx,2'bxx} : dec_ma_data_BCop12 = 1'b1;  /* MOV,word[BC],A */
                {8'h79,8'hxx,2'bxx} : dec_ma_data_BCop12 = 1'b1;  /* MOVW,AX,word[BC] */
                {8'h78,8'hxx,2'bxx} : dec_ma_data_BCop12 = 1'b1;  /* MOVW,word[BC],AX */
                default : dec_ma_data_BCop12 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ma_data_Bop12;
    reg    dec_ma_data_Bop12;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_ma_data_Bop12 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h19,8'hxx,2'bxx} : dec_ma_data_Bop12 = 1'b1;  /* MOV,word[B],#byte */
                {8'h09,8'hxx,2'bxx} : dec_ma_data_Bop12 = 1'b1;  /* MOV,A,word[B] */
                {8'h18,8'hxx,2'bxx} : dec_ma_data_Bop12 = 1'b1;  /* MOV,word[B],A */
                {8'h59,8'hxx,2'bxx} : dec_ma_data_Bop12 = 1'b1;  /* MOVW,AX,word[B] */
                {8'h58,8'hxx,2'bxx} : dec_ma_data_Bop12 = 1'b1;  /* MOVW,word[B],AX */
                default : dec_ma_data_Bop12 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ma_data_Cop12;
    reg    dec_ma_data_Cop12;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_ma_data_Cop12 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h38,8'hxx,2'bxx} : dec_ma_data_Cop12 = 1'b1;  /* MOV,word[C],#byte */
                {8'h29,8'hxx,2'bxx} : dec_ma_data_Cop12 = 1'b1;  /* MOV,A,word[C] */
                {8'h28,8'hxx,2'bxx} : dec_ma_data_Cop12 = 1'b1;  /* MOV,word[C],A */
                {8'h69,8'hxx,2'bxx} : dec_ma_data_Cop12 = 1'b1;  /* MOVW,AX,word[C] */
                {8'h68,8'hxx,2'bxx} : dec_ma_data_Cop12 = 1'b1;  /* MOVW,word[C],AX */
                default : dec_ma_data_Cop12 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_sp_set_enable;
    reg    dec_sp_set_enable;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(decout_mask == 1'b1) begin
//            dec_sp_set_enable = 1'b0;
//        end else if(rstvec == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1) begin
            dec_sp_set_enable = 1'b0;
        end else if(ivack == 1'b1) begin
            casex ({stage_adr})  
                {2'b00} : dec_sp_set_enable = 1'b1;  /* Interrupt */
                {2'b01} : dec_sp_set_enable = 1'b1;  /* Interrupt */
                default : dec_sp_set_enable = 1'b0;
            endcase
        end else if(skpack == 1'b1) begin
            dec_sp_set_enable = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hca,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALL,,AX */
                {8'h61,8'hca,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALL,,AX */
                {8'h61,8'hda,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALL,,BC */
                {8'h61,8'hda,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALL,,BC */
                {8'h61,8'hea,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALL,,DE */
                {8'h61,8'hea,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALL,,DE */
                {8'h61,8'hfa,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALL,,HL */
                {8'h61,8'hfa,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALL,,HL */
                {8'hfe,8'hxx,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALL,,$!addr16 */
                {8'hfe,8'hxx,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALL,,$!addr16 */
                {8'hfd,8'hxx,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALL,,!addr16 */
                {8'hfd,8'hxx,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALL,,!addr16 */
                {8'hfc,8'hxx,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALL,,!!addr20 */
                {8'hfc,8'hxx,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALL,,!!addr20 */
                {8'h61,8'h84,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[0080h] */
                {8'h61,8'h84,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[0080h] */
                {8'h61,8'h94,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[0082h] */
                {8'h61,8'h94,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[0082h] */
                {8'h61,8'ha4,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[0084h] */
                {8'h61,8'ha4,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[0084h] */
                {8'h61,8'hb4,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[0086h] */
                {8'h61,8'hb4,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[0086h] */
                {8'h61,8'hc4,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[0088h] */
                {8'h61,8'hc4,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[0088h] */
                {8'h61,8'hd4,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[008Ah] */
                {8'h61,8'hd4,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[008Ah] */
                {8'h61,8'he4,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[008Ch] */
                {8'h61,8'he4,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[008Ch] */
                {8'h61,8'hf4,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[008Eh] */
                {8'h61,8'hf4,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[008Eh] */
                {8'h61,8'h85,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[0090h] */
                {8'h61,8'h85,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[0090h] */
                {8'h61,8'h95,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[0092h] */
                {8'h61,8'h95,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[0092h] */
                {8'h61,8'ha5,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[0094h] */
                {8'h61,8'ha5,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[0094h] */
                {8'h61,8'hb5,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[0096h] */
                {8'h61,8'hb5,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[0096h] */
                {8'h61,8'hc5,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[0098h] */
                {8'h61,8'hc5,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[0098h] */
                {8'h61,8'hd5,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[009Ah] */
                {8'h61,8'hd5,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[009Ah] */
                {8'h61,8'he5,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[009Ch] */
                {8'h61,8'he5,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[009Ch] */
                {8'h61,8'hf5,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[009Eh] */
                {8'h61,8'hf5,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[009Eh] */
                {8'h61,8'h86,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00A0h] */
                {8'h61,8'h86,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00A0h] */
                {8'h61,8'h96,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00A2h] */
                {8'h61,8'h96,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00A2h] */
                {8'h61,8'ha6,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00A4h] */
                {8'h61,8'ha6,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00A4h] */
                {8'h61,8'hb6,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00A6h] */
                {8'h61,8'hb6,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00A6h] */
                {8'h61,8'hc6,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00A8h] */
                {8'h61,8'hc6,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00A8h] */
                {8'h61,8'hd6,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00AAh] */
                {8'h61,8'hd6,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00AAh] */
                {8'h61,8'he6,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00ACh] */
                {8'h61,8'he6,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00ACh] */
                {8'h61,8'hf6,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00AEh] */
                {8'h61,8'hf6,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00AEh] */
                {8'h61,8'h87,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00B0h] */
                {8'h61,8'h87,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00B0h] */
                {8'h61,8'h97,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00B2h] */
                {8'h61,8'h97,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00B2h] */
                {8'h61,8'ha7,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00B4h] */
                {8'h61,8'ha7,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00B4h] */
                {8'h61,8'hb7,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00B6h] */
                {8'h61,8'hb7,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00B6h] */
                {8'h61,8'hc7,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00B8h] */
                {8'h61,8'hc7,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00B8h] */
                {8'h61,8'hd7,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00BAh] */
                {8'h61,8'hd7,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00BAh] */
                {8'h61,8'he7,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00BCh] */
                {8'h61,8'he7,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00BCh] */
                {8'h61,8'hf7,2'bx0} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00BEh] */
                {8'h61,8'hf7,2'bx1} : dec_sp_set_enable = 1'b1;  /* CALLT,,[00BEh] */
                {8'h61,8'hcc,2'bx0} : dec_sp_set_enable = 1'b1;  /* BRK,, */
                {8'h61,8'hcc,2'bx1} : dec_sp_set_enable = 1'b1;  /* BRK,, */
                {8'hd7,8'hxx,2'b00} : dec_sp_set_enable = 1'b1;  /* RET,, */
                {8'hd7,8'hxx,2'b01} : dec_sp_set_enable = 1'b1;  /* RET,, */
                {8'h61,8'hec,2'b00} : dec_sp_set_enable = 1'b1;  /* RETB,, */
                {8'h61,8'hec,2'b01} : dec_sp_set_enable = 1'b1;  /* RETB,, */
                {8'h61,8'hfc,2'b00} : dec_sp_set_enable = 1'b1;  /* RETI,, */
                {8'h61,8'hfc,2'b01} : dec_sp_set_enable = 1'b1;  /* RETI,, */
                {8'h61,8'hdd,2'bxx} : dec_sp_set_enable = 1'b1;  /* PUSH,,PSW */
                {8'hc1,8'hxx,2'bxx} : dec_sp_set_enable = 1'b1;  /* PUSH,,AX */
                {8'hc3,8'hxx,2'bxx} : dec_sp_set_enable = 1'b1;  /* PUSH,,BC */
                {8'hc5,8'hxx,2'bxx} : dec_sp_set_enable = 1'b1;  /* PUSH,,DE */
                {8'hc7,8'hxx,2'bxx} : dec_sp_set_enable = 1'b1;  /* PUSH,,HL */
                {8'h61,8'hcd,2'bxx} : dec_sp_set_enable = 1'b1;  /* POP,,PSW */
                {8'hc0,8'hxx,2'bxx} : dec_sp_set_enable = 1'b1;  /* POP,,AX */
                {8'hc2,8'hxx,2'bxx} : dec_sp_set_enable = 1'b1;  /* POP,,BC */
                {8'hc4,8'hxx,2'bxx} : dec_sp_set_enable = 1'b1;  /* POP,,DE */
                {8'hc6,8'hxx,2'bxx} : dec_sp_set_enable = 1'b1;  /* POP,,HL */
                {8'hff,8'hxx,2'bx0} : dec_sp_set_enable = 1'b1;  /* SOFT,,BREAK */
                {8'hff,8'hxx,2'bx1} : dec_sp_set_enable = 1'b1;  /* SOFT,,BREAK */
                {8'h61,8'ha1,2'bx0} : dec_sp_set_enable = 1'b1;  /* SOFT2,,BREAK */
                {8'h61,8'ha1,2'bx1} : dec_sp_set_enable = 1'b1;  /* SOFT2,,BREAK */
                {8'h61,8'hb1,2'bx0} : dec_sp_set_enable = 1'b1;  /* SOFT3,,BREAK */
                {8'h61,8'hb1,2'bx1} : dec_sp_set_enable = 1'b1;  /* SOFT3,,BREAK */
                {8'h61,8'hc1,2'bx0} : dec_sp_set_enable = 1'b1;  /* SOFT4,,BREAK */
                {8'h61,8'hc1,2'bx1} : dec_sp_set_enable = 1'b1;  /* SOFT4,,BREAK */
                default : dec_sp_set_enable = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_sp_inc;
    reg    dec_sp_inc;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_sp_inc = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'hd7,8'hxx,2'b00} : dec_sp_inc = 1'b1;  /* RET,, */
                {8'hd7,8'hxx,2'b01} : dec_sp_inc = 1'b1;  /* RET,, */
                {8'h61,8'hec,2'b00} : dec_sp_inc = 1'b1;  /* RETB,, */
                {8'h61,8'hec,2'b01} : dec_sp_inc = 1'b1;  /* RETB,, */
                {8'h61,8'hfc,2'b00} : dec_sp_inc = 1'b1;  /* RETI,, */
                {8'h61,8'hfc,2'b01} : dec_sp_inc = 1'b1;  /* RETI,, */
                {8'h61,8'hcd,2'bxx} : dec_sp_inc = 1'b1;  /* POP,,PSW */
                {8'hc0,8'hxx,2'bxx} : dec_sp_inc = 1'b1;  /* POP,,AX */
                {8'hc2,8'hxx,2'bxx} : dec_sp_inc = 1'b1;  /* POP,,BC */
                {8'hc4,8'hxx,2'bxx} : dec_sp_inc = 1'b1;  /* POP,,DE */
                {8'hc6,8'hxx,2'bxx} : dec_sp_inc = 1'b1;  /* POP,,HL */
                default : dec_sp_inc = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_sp_dec;
    reg    dec_sp_dec;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(decout_mask == 1'b1) begin
//            dec_sp_dec = 1'b0;
//        end else if(rstvec == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1) begin
            dec_sp_dec = 1'b0;
        end else if(ivack == 1'b1) begin
            casex ({stage_adr})  
                {2'b00} : dec_sp_dec = 1'b1;  /* Interrupt */
                {2'b01} : dec_sp_dec = 1'b1;  /* Interrupt */
                default : dec_sp_dec = 1'b0;
            endcase
        end else if(skpack == 1'b1) begin
            dec_sp_dec = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hca,2'bx0} : dec_sp_dec = 1'b1;  /* CALL,,AX */
                {8'h61,8'hca,2'bx1} : dec_sp_dec = 1'b1;  /* CALL,,AX */
                {8'h61,8'hda,2'bx0} : dec_sp_dec = 1'b1;  /* CALL,,BC */
                {8'h61,8'hda,2'bx1} : dec_sp_dec = 1'b1;  /* CALL,,BC */
                {8'h61,8'hea,2'bx0} : dec_sp_dec = 1'b1;  /* CALL,,DE */
                {8'h61,8'hea,2'bx1} : dec_sp_dec = 1'b1;  /* CALL,,DE */
                {8'h61,8'hfa,2'bx0} : dec_sp_dec = 1'b1;  /* CALL,,HL */
                {8'h61,8'hfa,2'bx1} : dec_sp_dec = 1'b1;  /* CALL,,HL */
                {8'hfe,8'hxx,2'bx0} : dec_sp_dec = 1'b1;  /* CALL,,$!addr16 */
                {8'hfe,8'hxx,2'bx1} : dec_sp_dec = 1'b1;  /* CALL,,$!addr16 */
                {8'hfd,8'hxx,2'bx0} : dec_sp_dec = 1'b1;  /* CALL,,!addr16 */
                {8'hfd,8'hxx,2'bx1} : dec_sp_dec = 1'b1;  /* CALL,,!addr16 */
                {8'hfc,8'hxx,2'bx0} : dec_sp_dec = 1'b1;  /* CALL,,!!addr20 */
                {8'hfc,8'hxx,2'bx1} : dec_sp_dec = 1'b1;  /* CALL,,!!addr20 */
                {8'h61,8'h84,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[0080h] */
                {8'h61,8'h84,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[0080h] */
                {8'h61,8'h94,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[0082h] */
                {8'h61,8'h94,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[0082h] */
                {8'h61,8'ha4,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[0084h] */
                {8'h61,8'ha4,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[0084h] */
                {8'h61,8'hb4,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[0086h] */
                {8'h61,8'hb4,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[0086h] */
                {8'h61,8'hc4,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[0088h] */
                {8'h61,8'hc4,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[0088h] */
                {8'h61,8'hd4,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[008Ah] */
                {8'h61,8'hd4,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[008Ah] */
                {8'h61,8'he4,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[008Ch] */
                {8'h61,8'he4,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[008Ch] */
                {8'h61,8'hf4,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[008Eh] */
                {8'h61,8'hf4,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[008Eh] */
                {8'h61,8'h85,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[0090h] */
                {8'h61,8'h85,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[0090h] */
                {8'h61,8'h95,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[0092h] */
                {8'h61,8'h95,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[0092h] */
                {8'h61,8'ha5,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[0094h] */
                {8'h61,8'ha5,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[0094h] */
                {8'h61,8'hb5,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[0096h] */
                {8'h61,8'hb5,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[0096h] */
                {8'h61,8'hc5,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[0098h] */
                {8'h61,8'hc5,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[0098h] */
                {8'h61,8'hd5,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[009Ah] */
                {8'h61,8'hd5,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[009Ah] */
                {8'h61,8'he5,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[009Ch] */
                {8'h61,8'he5,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[009Ch] */
                {8'h61,8'hf5,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[009Eh] */
                {8'h61,8'hf5,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[009Eh] */
                {8'h61,8'h86,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[00A0h] */
                {8'h61,8'h86,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[00A0h] */
                {8'h61,8'h96,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[00A2h] */
                {8'h61,8'h96,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[00A2h] */
                {8'h61,8'ha6,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[00A4h] */
                {8'h61,8'ha6,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[00A4h] */
                {8'h61,8'hb6,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[00A6h] */
                {8'h61,8'hb6,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[00A6h] */
                {8'h61,8'hc6,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[00A8h] */
                {8'h61,8'hc6,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[00A8h] */
                {8'h61,8'hd6,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[00AAh] */
                {8'h61,8'hd6,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[00AAh] */
                {8'h61,8'he6,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[00ACh] */
                {8'h61,8'he6,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[00ACh] */
                {8'h61,8'hf6,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[00AEh] */
                {8'h61,8'hf6,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[00AEh] */
                {8'h61,8'h87,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[00B0h] */
                {8'h61,8'h87,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[00B0h] */
                {8'h61,8'h97,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[00B2h] */
                {8'h61,8'h97,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[00B2h] */
                {8'h61,8'ha7,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[00B4h] */
                {8'h61,8'ha7,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[00B4h] */
                {8'h61,8'hb7,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[00B6h] */
                {8'h61,8'hb7,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[00B6h] */
                {8'h61,8'hc7,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[00B8h] */
                {8'h61,8'hc7,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[00B8h] */
                {8'h61,8'hd7,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[00BAh] */
                {8'h61,8'hd7,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[00BAh] */
                {8'h61,8'he7,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[00BCh] */
                {8'h61,8'he7,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[00BCh] */
                {8'h61,8'hf7,2'bx0} : dec_sp_dec = 1'b1;  /* CALLT,,[00BEh] */
                {8'h61,8'hf7,2'bx1} : dec_sp_dec = 1'b1;  /* CALLT,,[00BEh] */
                {8'h61,8'hcc,2'bx0} : dec_sp_dec = 1'b1;  /* BRK,, */
                {8'h61,8'hcc,2'bx1} : dec_sp_dec = 1'b1;  /* BRK,, */
                {8'h61,8'hdd,2'bxx} : dec_sp_dec = 1'b1;  /* PUSH,,PSW */
                {8'hc1,8'hxx,2'bxx} : dec_sp_dec = 1'b1;  /* PUSH,,AX */
                {8'hc3,8'hxx,2'bxx} : dec_sp_dec = 1'b1;  /* PUSH,,BC */
                {8'hc5,8'hxx,2'bxx} : dec_sp_dec = 1'b1;  /* PUSH,,DE */
                {8'hc7,8'hxx,2'bxx} : dec_sp_dec = 1'b1;  /* PUSH,,HL */
                {8'hff,8'hxx,2'bx0} : dec_sp_dec = 1'b1;  /* SOFT,,BREAK */
                {8'hff,8'hxx,2'bx1} : dec_sp_dec = 1'b1;  /* SOFT,,BREAK */
                {8'h61,8'ha1,2'bx0} : dec_sp_dec = 1'b1;  /* SOFT2,,BREAK */
                {8'h61,8'ha1,2'bx1} : dec_sp_dec = 1'b1;  /* SOFT2,,BREAK */
                {8'h61,8'hb1,2'bx0} : dec_sp_dec = 1'b1;  /* SOFT3,,BREAK */
                {8'h61,8'hb1,2'bx1} : dec_sp_dec = 1'b1;  /* SOFT3,,BREAK */
                {8'h61,8'hc1,2'bx0} : dec_sp_dec = 1'b1;  /* SOFT4,,BREAK */
                {8'h61,8'hc1,2'bx1} : dec_sp_dec = 1'b1;  /* SOFT4,,BREAK */
                default : dec_sp_dec = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_pc_inc1;
    reg    dec_pc_inc1;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1) begin
            dec_pc_inc1 = 1'b0;
        end else if(skpack == 1'b1) begin
            casex ({ID_stage0,ID_stage1})  
                {8'h60,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOV,A,X */
                {8'h62,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOV,A,C */
                {8'h63,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOV,A,B */
                {8'h64,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOV,A,E */
                {8'h65,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOV,A,D */
                {8'h66,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOV,A,L */
                {8'h67,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOV,A,H */
                {8'h70,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOV,X,A */
                {8'h72,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOV,C,A */
                {8'h73,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOV,B,A */
                {8'h74,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOV,E,A */
                {8'h75,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOV,D,A */
                {8'h76,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOV,L,A */
                {8'h77,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOV,H,A */
                {8'h89,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOV,A,[DE] */
                {8'h99,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOV,[DE],A */
                {8'h8b,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOV,A,[HL] */
                {8'h9b,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOV,[HL],A */
                {8'h08,8'hxx} : dec_pc_inc1 = 1'b1;  /* XCH,A,X */
                {8'he1,8'hxx} : dec_pc_inc1 = 1'b1;  /* ONEB,,A */
                {8'he0,8'hxx} : dec_pc_inc1 = 1'b1;  /* ONEB,,X */
                {8'he3,8'hxx} : dec_pc_inc1 = 1'b1;  /* ONEB,,B */
                {8'he2,8'hxx} : dec_pc_inc1 = 1'b1;  /* ONEB,,C */
                {8'hf1,8'hxx} : dec_pc_inc1 = 1'b1;  /* CLRB,,A */
                {8'hf0,8'hxx} : dec_pc_inc1 = 1'b1;  /* CLRB,,X */
                {8'hf3,8'hxx} : dec_pc_inc1 = 1'b1;  /* CLRB,,B */
                {8'hf2,8'hxx} : dec_pc_inc1 = 1'b1;  /* CLRB,,C */
                {8'h13,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOVW,AX,BC */
                {8'h12,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOVW,BC,AX */
                {8'h15,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOVW,AX,DE */
                {8'h14,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOVW,DE,AX */
                {8'h17,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOVW,AX,HL */
                {8'h16,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOVW,HL,AX */
                {8'ha9,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOVW,AX,[DE] */
                {8'hb9,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOVW,[DE],AX */
                {8'hab,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOVW,AX,[HL] */
                {8'hbb,8'hxx} : dec_pc_inc1 = 1'b1;  /* MOVW,[HL],AX */
                {8'h33,8'hxx} : dec_pc_inc1 = 1'b1;  /* XCHW,AX,BC */
                {8'h35,8'hxx} : dec_pc_inc1 = 1'b1;  /* XCHW,AX,DE */
                {8'h37,8'hxx} : dec_pc_inc1 = 1'b1;  /* XCHW,AX,HL */
                {8'he6,8'hxx} : dec_pc_inc1 = 1'b1;  /* ONEW,,AX */
                {8'he7,8'hxx} : dec_pc_inc1 = 1'b1;  /* ONEW,,BC */
                {8'hf6,8'hxx} : dec_pc_inc1 = 1'b1;  /* CLRW,,AX */
                {8'hf7,8'hxx} : dec_pc_inc1 = 1'b1;  /* CLRW,,BC */
                {8'h0d,8'hxx} : dec_pc_inc1 = 1'b1;  /* ADD,A,[HL] */
                {8'h1d,8'hxx} : dec_pc_inc1 = 1'b1;  /* ADDC,A,[HL] */
                {8'h2d,8'hxx} : dec_pc_inc1 = 1'b1;  /* SUB,A,[HL] */
                {8'h3d,8'hxx} : dec_pc_inc1 = 1'b1;  /* SUBC,A,[HL] */
                {8'h5d,8'hxx} : dec_pc_inc1 = 1'b1;  /* AND,A,[HL] */
                {8'h6d,8'hxx} : dec_pc_inc1 = 1'b1;  /* OR,A,[HL] */
                {8'h7d,8'hxx} : dec_pc_inc1 = 1'b1;  /* XOR,A,[HL] */
                {8'h4d,8'hxx} : dec_pc_inc1 = 1'b1;  /* CMP,A,[HL] */
                {8'hd1,8'hxx} : dec_pc_inc1 = 1'b1;  /* CMP0,,A */
                {8'hd0,8'hxx} : dec_pc_inc1 = 1'b1;  /* CMP0,,X */
                {8'hd3,8'hxx} : dec_pc_inc1 = 1'b1;  /* CMP0,,B */
                {8'hd2,8'hxx} : dec_pc_inc1 = 1'b1;  /* CMP0,,C */
                {8'h01,8'hxx} : dec_pc_inc1 = 1'b1;  /* ADDW,AX,AX */
                {8'h03,8'hxx} : dec_pc_inc1 = 1'b1;  /* ADDW,AX,BC */
                {8'h05,8'hxx} : dec_pc_inc1 = 1'b1;  /* ADDW,AX,DE */
                {8'h07,8'hxx} : dec_pc_inc1 = 1'b1;  /* ADDW,AX,HL */
                {8'h21,8'hxx} : dec_pc_inc1 = 1'b1;  /* SUBW,AX,AX */
                {8'h23,8'hxx} : dec_pc_inc1 = 1'b1;  /* SUBW,AX,BC */
                {8'h25,8'hxx} : dec_pc_inc1 = 1'b1;  /* SUBW,AX,DE */
                {8'h27,8'hxx} : dec_pc_inc1 = 1'b1;  /* SUBW,AX,HL */
                {8'h43,8'hxx} : dec_pc_inc1 = 1'b1;  /* CMPW,AX,BC */
                {8'h45,8'hxx} : dec_pc_inc1 = 1'b1;  /* CMPW,AX,DE */
                {8'h47,8'hxx} : dec_pc_inc1 = 1'b1;  /* CMPW,AX,HL */
                {8'hd6,8'hxx} : dec_pc_inc1 = 1'b1;  /* MULU,,X */
                {8'h80,8'hxx} : dec_pc_inc1 = 1'b1;  /* INC,,X */
                {8'h81,8'hxx} : dec_pc_inc1 = 1'b1;  /* INC,,A */
                {8'h82,8'hxx} : dec_pc_inc1 = 1'b1;  /* INC,,C */
                {8'h83,8'hxx} : dec_pc_inc1 = 1'b1;  /* INC,,B */
                {8'h84,8'hxx} : dec_pc_inc1 = 1'b1;  /* INC,,E */
                {8'h85,8'hxx} : dec_pc_inc1 = 1'b1;  /* INC,,D */
                {8'h86,8'hxx} : dec_pc_inc1 = 1'b1;  /* INC,,L */
                {8'h87,8'hxx} : dec_pc_inc1 = 1'b1;  /* INC,,H */
                {8'h90,8'hxx} : dec_pc_inc1 = 1'b1;  /* DEC,,X */
                {8'h91,8'hxx} : dec_pc_inc1 = 1'b1;  /* DEC,,A */
                {8'h92,8'hxx} : dec_pc_inc1 = 1'b1;  /* DEC,,C */
                {8'h93,8'hxx} : dec_pc_inc1 = 1'b1;  /* DEC,,B */
                {8'h94,8'hxx} : dec_pc_inc1 = 1'b1;  /* DEC,,E */
                {8'h95,8'hxx} : dec_pc_inc1 = 1'b1;  /* DEC,,D */
                {8'h96,8'hxx} : dec_pc_inc1 = 1'b1;  /* DEC,,L */
                {8'h97,8'hxx} : dec_pc_inc1 = 1'b1;  /* DEC,,H */
                {8'ha1,8'hxx} : dec_pc_inc1 = 1'b1;  /* INCW,,AX */
                {8'ha3,8'hxx} : dec_pc_inc1 = 1'b1;  /* INCW,,BC */
                {8'ha5,8'hxx} : dec_pc_inc1 = 1'b1;  /* INCW,,DE */
                {8'ha7,8'hxx} : dec_pc_inc1 = 1'b1;  /* INCW,,HL */
                {8'hb1,8'hxx} : dec_pc_inc1 = 1'b1;  /* DECW,,AX */
                {8'hb3,8'hxx} : dec_pc_inc1 = 1'b1;  /* DECW,,BC */
                {8'hb5,8'hxx} : dec_pc_inc1 = 1'b1;  /* DECW,,DE */
                {8'hb7,8'hxx} : dec_pc_inc1 = 1'b1;  /* DECW,,HL */
                {8'hd7,8'hxx} : dec_pc_inc1 = 1'b1;  /* RET,, */
                {8'hc1,8'hxx} : dec_pc_inc1 = 1'b1;  /* PUSH,,AX */
                {8'hc3,8'hxx} : dec_pc_inc1 = 1'b1;  /* PUSH,,BC */
                {8'hc5,8'hxx} : dec_pc_inc1 = 1'b1;  /* PUSH,,DE */
                {8'hc7,8'hxx} : dec_pc_inc1 = 1'b1;  /* PUSH,,HL */
                {8'hc0,8'hxx} : dec_pc_inc1 = 1'b1;  /* POP,,AX */
                {8'hc2,8'hxx} : dec_pc_inc1 = 1'b1;  /* POP,,BC */
                {8'hc4,8'hxx} : dec_pc_inc1 = 1'b1;  /* POP,,DE */
                {8'hc6,8'hxx} : dec_pc_inc1 = 1'b1;  /* POP,,HL */
                {8'h00,8'hxx} : dec_pc_inc1 = 1'b1;  /* NOP,, */
                {8'h11,8'hxx} : dec_pc_inc1 = 1'b1;  /* PREFIX,, */
                {8'hff,8'hxx} : dec_pc_inc1 = 1'b1;  /* SOFT,,BREAK */
                default : dec_pc_inc1 = 1'b0;
            endcase
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h60,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOV,A,X */
                {8'h62,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOV,A,C */
                {8'h63,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOV,A,B */
                {8'h64,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOV,A,E */
                {8'h65,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOV,A,D */
                {8'h66,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOV,A,L */
                {8'h67,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOV,A,H */
                {8'h70,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOV,X,A */
                {8'h72,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOV,C,A */
                {8'h73,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOV,B,A */
                {8'h74,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOV,E,A */
                {8'h75,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOV,D,A */
                {8'h76,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOV,L,A */
                {8'h77,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOV,H,A */
                {8'h89,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOV,A,[DE] */
                {8'h99,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOV,[DE],A */
                {8'h8b,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOV,A,[HL] */
                {8'h9b,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOV,[HL],A */
                {8'h08,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* XCH,A,X */
                {8'he1,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* ONEB,,A */
                {8'he0,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* ONEB,,X */
                {8'he3,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* ONEB,,B */
                {8'he2,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* ONEB,,C */
                {8'hf1,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* CLRB,,A */
                {8'hf0,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* CLRB,,X */
                {8'hf3,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* CLRB,,B */
                {8'hf2,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* CLRB,,C */
                {8'h13,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOVW,AX,BC */
                {8'h12,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOVW,BC,AX */
                {8'h15,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOVW,AX,DE */
                {8'h14,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOVW,DE,AX */
                {8'h17,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOVW,AX,HL */
                {8'h16,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOVW,HL,AX */
                {8'ha9,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOVW,AX,[DE] */
                {8'hb9,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOVW,[DE],AX */
                {8'hab,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOVW,AX,[HL] */
                {8'hbb,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MOVW,[HL],AX */
                {8'h33,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* XCHW,AX,BC */
                {8'h35,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* XCHW,AX,DE */
                {8'h37,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* XCHW,AX,HL */
                {8'he6,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* ONEW,,AX */
                {8'he7,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* ONEW,,BC */
                {8'hf6,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* CLRW,,AX */
                {8'hf7,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* CLRW,,BC */
                {8'h0d,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* ADD,A,[HL] */
                {8'h1d,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* ADDC,A,[HL] */
                {8'h2d,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* SUB,A,[HL] */
                {8'h3d,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* SUBC,A,[HL] */
                {8'h5d,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* AND,A,[HL] */
                {8'h6d,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* OR,A,[HL] */
                {8'h7d,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* XOR,A,[HL] */
                {8'h4d,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* CMP,A,[HL] */
                {8'hd1,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* CMP0,,A */
                {8'hd0,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* CMP0,,X */
                {8'hd3,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* CMP0,,B */
                {8'hd2,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* CMP0,,C */
                {8'h01,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* ADDW,AX,AX */
                {8'h03,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* ADDW,AX,BC */
                {8'h05,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* ADDW,AX,DE */
                {8'h07,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* ADDW,AX,HL */
                {8'h21,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* SUBW,AX,AX */
                {8'h23,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* SUBW,AX,BC */
                {8'h25,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* SUBW,AX,DE */
                {8'h27,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* SUBW,AX,HL */
                {8'h43,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* CMPW,AX,BC */
                {8'h45,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* CMPW,AX,DE */
                {8'h47,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* CMPW,AX,HL */
                {8'hd6,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* MULU,,X */
                {8'h80,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* INC,,X */
                {8'h81,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* INC,,A */
                {8'h82,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* INC,,C */
                {8'h83,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* INC,,B */
                {8'h84,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* INC,,E */
                {8'h85,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* INC,,D */
                {8'h86,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* INC,,L */
                {8'h87,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* INC,,H */
                {8'h90,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* DEC,,X */
                {8'h91,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* DEC,,A */
                {8'h92,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* DEC,,C */
                {8'h93,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* DEC,,B */
                {8'h94,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* DEC,,E */
                {8'h95,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* DEC,,D */
                {8'h96,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* DEC,,L */
                {8'h97,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* DEC,,H */
                {8'ha1,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* INCW,,AX */
                {8'ha3,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* INCW,,BC */
                {8'ha5,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* INCW,,DE */
                {8'ha7,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* INCW,,HL */
                {8'hb1,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* DECW,,AX */
                {8'hb3,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* DECW,,BC */
                {8'hb5,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* DECW,,DE */
                {8'hb7,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* DECW,,HL */
                {8'hc1,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* PUSH,,AX */
                {8'hc3,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* PUSH,,BC */
                {8'hc5,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* PUSH,,DE */
                {8'hc7,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* PUSH,,HL */
                {8'hc0,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* POP,,AX */
                {8'hc2,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* POP,,BC */
                {8'hc4,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* POP,,DE */
                {8'hc6,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* POP,,HL */
                {8'h00,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* NOP,, */
                {8'h11,8'hxx,2'bxx} : dec_pc_inc1 = 1'b1;  /* PREFIX,, */
                {8'hff,8'hxx,2'bx0} : dec_pc_inc1 = 1'b1;  /* SOFT,,BREAK */
                default : dec_pc_inc1 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_pc_inc2;
    reg    dec_pc_inc2;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1) begin
            dec_pc_inc2 = 1'b0;
        end else if(skpack == 1'b1) begin
            casex ({ID_stage0,ID_stage1})  
                {8'h50,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOV,X,#byte */
                {8'h51,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOV,A,#byte */
                {8'h52,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOV,C,#byte */
                {8'h53,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOV,B,#byte */
                {8'h54,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOV,E,#byte */
                {8'h55,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOV,D,#byte */
                {8'h56,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOV,L,#byte */
                {8'h57,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOV,H,#byte */
                {8'h8d,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOV,A,saddr */
                {8'h9d,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOV,saddr,A */
                {8'h8e,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOV,A,sfr */
                {8'h9e,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOV,sfr,A */
                {8'h41,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOV,ES,#byte */
                {8'h8a,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOV,A,[DE+byte] */
                {8'h9a,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOV,[DE+byte],A */
                {8'h8c,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOV,A,[HL+byte] */
                {8'h9c,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOV,[HL+byte],A */
                {8'h61,8'hc9} : dec_pc_inc2 = 1'b1;  /* MOV,A,[HL+B] */
                {8'h61,8'hd9} : dec_pc_inc2 = 1'b1;  /* MOV,[HL+B],A */
                {8'h61,8'he9} : dec_pc_inc2 = 1'b1;  /* MOV,A,[HL+C] */
                {8'h61,8'hf9} : dec_pc_inc2 = 1'b1;  /* MOV,[HL+C],A */
                {8'h88,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOV,A,[SP+byte] */
                {8'h98,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOV,[SP+byte],A */
                {8'he8,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOV,B,saddr */
                {8'hf8,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOV,C,saddr */
                {8'hd8,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOV,X,saddr */
                {8'h61,8'h8a} : dec_pc_inc2 = 1'b1;  /* XCH,A,C */
                {8'h61,8'h8b} : dec_pc_inc2 = 1'b1;  /* XCH,A,B */
                {8'h61,8'h8c} : dec_pc_inc2 = 1'b1;  /* XCH,A,E */
                {8'h61,8'h8d} : dec_pc_inc2 = 1'b1;  /* XCH,A,D */
                {8'h61,8'h8e} : dec_pc_inc2 = 1'b1;  /* XCH,A,L */
                {8'h61,8'h8f} : dec_pc_inc2 = 1'b1;  /* XCH,A,H */
                {8'h61,8'hae} : dec_pc_inc2 = 1'b1;  /* XCH,A,[DE] */
                {8'h61,8'hac} : dec_pc_inc2 = 1'b1;  /* XCH,A,[HL] */
                {8'h61,8'hb9} : dec_pc_inc2 = 1'b1;  /* XCH,A,[HL+B] */
                {8'h61,8'ha9} : dec_pc_inc2 = 1'b1;  /* XCH,A,[HL+C] */
                {8'he4,8'hxx} : dec_pc_inc2 = 1'b1;  /* ONEB,,saddr */
                {8'hf4,8'hxx} : dec_pc_inc2 = 1'b1;  /* CLRB,,saddr */
                {8'had,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOVW,AX,saddrp */
                {8'hbd,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOVW,saddrp,AX */
                {8'hae,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOVW,AX,sfrp */
                {8'hbe,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOVW,sfrp,AX */
                {8'haa,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOVW,AX,[DE+byte] */
                {8'hba,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOVW,[DE+byte],AX */
                {8'hac,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOVW,AX,[HL+byte] */
                {8'hbc,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOVW,[HL+byte],AX */
                {8'ha8,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOVW,AX,[SP+byte] */
                {8'hb8,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOVW,[SP+byte],AX */
                {8'hda,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOVW,BC,saddrp */
                {8'hea,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOVW,DE,saddrp */
                {8'hfa,8'hxx} : dec_pc_inc2 = 1'b1;  /* MOVW,HL,saddrp */
                {8'h0c,8'hxx} : dec_pc_inc2 = 1'b1;  /* ADD,A,#byte */
                {8'h61,8'h08} : dec_pc_inc2 = 1'b1;  /* ADD,A,X */
                {8'h61,8'h0a} : dec_pc_inc2 = 1'b1;  /* ADD,A,C */
                {8'h61,8'h0b} : dec_pc_inc2 = 1'b1;  /* ADD,A,B */
                {8'h61,8'h0c} : dec_pc_inc2 = 1'b1;  /* ADD,A,E */
                {8'h61,8'h0d} : dec_pc_inc2 = 1'b1;  /* ADD,A,D */
                {8'h61,8'h0e} : dec_pc_inc2 = 1'b1;  /* ADD,A,L */
                {8'h61,8'h0f} : dec_pc_inc2 = 1'b1;  /* ADD,A,H */
                {8'h61,8'h00} : dec_pc_inc2 = 1'b1;  /* ADD,X,A */
                {8'h61,8'h01} : dec_pc_inc2 = 1'b1;  /* ADD,A,A */
                {8'h61,8'h02} : dec_pc_inc2 = 1'b1;  /* ADD,C,A */
                {8'h61,8'h03} : dec_pc_inc2 = 1'b1;  /* ADD,B,A */
                {8'h61,8'h04} : dec_pc_inc2 = 1'b1;  /* ADD,E,A */
                {8'h61,8'h05} : dec_pc_inc2 = 1'b1;  /* ADD,D,A */
                {8'h61,8'h06} : dec_pc_inc2 = 1'b1;  /* ADD,L,A */
                {8'h61,8'h07} : dec_pc_inc2 = 1'b1;  /* ADD,H,A */
                {8'h0b,8'hxx} : dec_pc_inc2 = 1'b1;  /* ADD,A,saddr */
                {8'h0e,8'hxx} : dec_pc_inc2 = 1'b1;  /* ADD,A,[HL+byte] */
                {8'h61,8'h80} : dec_pc_inc2 = 1'b1;  /* ADD,A,[HL+B] */
                {8'h61,8'h82} : dec_pc_inc2 = 1'b1;  /* ADD,A,[HL+C] */
                {8'h1c,8'hxx} : dec_pc_inc2 = 1'b1;  /* ADDC,A,#byte */
                {8'h61,8'h18} : dec_pc_inc2 = 1'b1;  /* ADDC,A,X */
                {8'h61,8'h1a} : dec_pc_inc2 = 1'b1;  /* ADDC,A,C */
                {8'h61,8'h1b} : dec_pc_inc2 = 1'b1;  /* ADDC,A,B */
                {8'h61,8'h1c} : dec_pc_inc2 = 1'b1;  /* ADDC,A,E */
                {8'h61,8'h1d} : dec_pc_inc2 = 1'b1;  /* ADDC,A,D */
                {8'h61,8'h1e} : dec_pc_inc2 = 1'b1;  /* ADDC,A,L */
                {8'h61,8'h1f} : dec_pc_inc2 = 1'b1;  /* ADDC,A,H */
                {8'h61,8'h10} : dec_pc_inc2 = 1'b1;  /* ADDC,X,A */
                {8'h61,8'h11} : dec_pc_inc2 = 1'b1;  /* ADDC,A,A */
                {8'h61,8'h12} : dec_pc_inc2 = 1'b1;  /* ADDC,C,A */
                {8'h61,8'h13} : dec_pc_inc2 = 1'b1;  /* ADDC,B,A */
                {8'h61,8'h14} : dec_pc_inc2 = 1'b1;  /* ADDC,E,A */
                {8'h61,8'h15} : dec_pc_inc2 = 1'b1;  /* ADDC,D,A */
                {8'h61,8'h16} : dec_pc_inc2 = 1'b1;  /* ADDC,L,A */
                {8'h61,8'h17} : dec_pc_inc2 = 1'b1;  /* ADDC,H,A */
                {8'h1b,8'hxx} : dec_pc_inc2 = 1'b1;  /* ADDC,A,saddr */
                {8'h1e,8'hxx} : dec_pc_inc2 = 1'b1;  /* ADDC,A,[HL+byte] */
                {8'h61,8'h90} : dec_pc_inc2 = 1'b1;  /* ADDC,A,[HL+B] */
                {8'h61,8'h92} : dec_pc_inc2 = 1'b1;  /* ADDC,A,[HL+C] */
                {8'h2c,8'hxx} : dec_pc_inc2 = 1'b1;  /* SUB,A,#byte */
                {8'h61,8'h28} : dec_pc_inc2 = 1'b1;  /* SUB,A,X */
                {8'h61,8'h2a} : dec_pc_inc2 = 1'b1;  /* SUB,A,C */
                {8'h61,8'h2b} : dec_pc_inc2 = 1'b1;  /* SUB,A,B */
                {8'h61,8'h2c} : dec_pc_inc2 = 1'b1;  /* SUB,A,E */
                {8'h61,8'h2d} : dec_pc_inc2 = 1'b1;  /* SUB,A,D */
                {8'h61,8'h2e} : dec_pc_inc2 = 1'b1;  /* SUB,A,L */
                {8'h61,8'h2f} : dec_pc_inc2 = 1'b1;  /* SUB,A,H */
                {8'h61,8'h20} : dec_pc_inc2 = 1'b1;  /* SUB,X,A */
                {8'h61,8'h21} : dec_pc_inc2 = 1'b1;  /* SUB,A,A */
                {8'h61,8'h22} : dec_pc_inc2 = 1'b1;  /* SUB,C,A */
                {8'h61,8'h23} : dec_pc_inc2 = 1'b1;  /* SUB,B,A */
                {8'h61,8'h24} : dec_pc_inc2 = 1'b1;  /* SUB,E,A */
                {8'h61,8'h25} : dec_pc_inc2 = 1'b1;  /* SUB,D,A */
                {8'h61,8'h26} : dec_pc_inc2 = 1'b1;  /* SUB,L,A */
                {8'h61,8'h27} : dec_pc_inc2 = 1'b1;  /* SUB,H,A */
                {8'h2b,8'hxx} : dec_pc_inc2 = 1'b1;  /* SUB,A,saddr */
                {8'h2e,8'hxx} : dec_pc_inc2 = 1'b1;  /* SUB,A,[HL+byte] */
                {8'h61,8'ha0} : dec_pc_inc2 = 1'b1;  /* SUB,A,[HL+B] */
                {8'h61,8'ha2} : dec_pc_inc2 = 1'b1;  /* SUB,A,[HL+C] */
                {8'h3c,8'hxx} : dec_pc_inc2 = 1'b1;  /* SUBC,A,#byte */
                {8'h61,8'h38} : dec_pc_inc2 = 1'b1;  /* SUBC,A,X */
                {8'h61,8'h3a} : dec_pc_inc2 = 1'b1;  /* SUBC,A,C */
                {8'h61,8'h3b} : dec_pc_inc2 = 1'b1;  /* SUBC,A,B */
                {8'h61,8'h3c} : dec_pc_inc2 = 1'b1;  /* SUBC,A,E */
                {8'h61,8'h3d} : dec_pc_inc2 = 1'b1;  /* SUBC,A,D */
                {8'h61,8'h3e} : dec_pc_inc2 = 1'b1;  /* SUBC,A,L */
                {8'h61,8'h3f} : dec_pc_inc2 = 1'b1;  /* SUBC,A,H */
                {8'h61,8'h30} : dec_pc_inc2 = 1'b1;  /* SUBC,X,A */
                {8'h61,8'h31} : dec_pc_inc2 = 1'b1;  /* SUBC,A,A */
                {8'h61,8'h32} : dec_pc_inc2 = 1'b1;  /* SUBC,C,A */
                {8'h61,8'h33} : dec_pc_inc2 = 1'b1;  /* SUBC,B,A */
                {8'h61,8'h34} : dec_pc_inc2 = 1'b1;  /* SUBC,E,A */
                {8'h61,8'h35} : dec_pc_inc2 = 1'b1;  /* SUBC,D,A */
                {8'h61,8'h36} : dec_pc_inc2 = 1'b1;  /* SUBC,L,A */
                {8'h61,8'h37} : dec_pc_inc2 = 1'b1;  /* SUBC,H,A */
                {8'h3b,8'hxx} : dec_pc_inc2 = 1'b1;  /* SUBC,A,saddr */
                {8'h3e,8'hxx} : dec_pc_inc2 = 1'b1;  /* SUBC,A,[HL+byte] */
                {8'h61,8'hb0} : dec_pc_inc2 = 1'b1;  /* SUBC,A,[HL+B] */
                {8'h61,8'hb2} : dec_pc_inc2 = 1'b1;  /* SUBC,A,[HL+C] */
                {8'h5c,8'hxx} : dec_pc_inc2 = 1'b1;  /* AND,A,#byte */
                {8'h61,8'h58} : dec_pc_inc2 = 1'b1;  /* AND,A,X */
                {8'h61,8'h5a} : dec_pc_inc2 = 1'b1;  /* AND,A,C */
                {8'h61,8'h5b} : dec_pc_inc2 = 1'b1;  /* AND,A,B */
                {8'h61,8'h5c} : dec_pc_inc2 = 1'b1;  /* AND,A,E */
                {8'h61,8'h5d} : dec_pc_inc2 = 1'b1;  /* AND,A,D */
                {8'h61,8'h5e} : dec_pc_inc2 = 1'b1;  /* AND,A,L */
                {8'h61,8'h5f} : dec_pc_inc2 = 1'b1;  /* AND,A,H */
                {8'h61,8'h50} : dec_pc_inc2 = 1'b1;  /* AND,X,A */
                {8'h61,8'h51} : dec_pc_inc2 = 1'b1;  /* AND,A,A */
                {8'h61,8'h52} : dec_pc_inc2 = 1'b1;  /* AND,C,A */
                {8'h61,8'h53} : dec_pc_inc2 = 1'b1;  /* AND,B,A */
                {8'h61,8'h54} : dec_pc_inc2 = 1'b1;  /* AND,E,A */
                {8'h61,8'h55} : dec_pc_inc2 = 1'b1;  /* AND,D,A */
                {8'h61,8'h56} : dec_pc_inc2 = 1'b1;  /* AND,L,A */
                {8'h61,8'h57} : dec_pc_inc2 = 1'b1;  /* AND,H,A */
                {8'h5b,8'hxx} : dec_pc_inc2 = 1'b1;  /* AND,A,saddr */
                {8'h5e,8'hxx} : dec_pc_inc2 = 1'b1;  /* AND,A,[HL+byte] */
                {8'h61,8'hd0} : dec_pc_inc2 = 1'b1;  /* AND,A,[HL+B] */
                {8'h61,8'hd2} : dec_pc_inc2 = 1'b1;  /* AND,A,[HL+C] */
                {8'h6c,8'hxx} : dec_pc_inc2 = 1'b1;  /* OR,A,#byte */
                {8'h61,8'h68} : dec_pc_inc2 = 1'b1;  /* OR,A,X */
                {8'h61,8'h6a} : dec_pc_inc2 = 1'b1;  /* OR,A,C */
                {8'h61,8'h6b} : dec_pc_inc2 = 1'b1;  /* OR,A,B */
                {8'h61,8'h6c} : dec_pc_inc2 = 1'b1;  /* OR,A,E */
                {8'h61,8'h6d} : dec_pc_inc2 = 1'b1;  /* OR,A,D */
                {8'h61,8'h6e} : dec_pc_inc2 = 1'b1;  /* OR,A,L */
                {8'h61,8'h6f} : dec_pc_inc2 = 1'b1;  /* OR,A,H */
                {8'h61,8'h60} : dec_pc_inc2 = 1'b1;  /* OR,X,A */
                {8'h61,8'h61} : dec_pc_inc2 = 1'b1;  /* OR,A,A */
                {8'h61,8'h62} : dec_pc_inc2 = 1'b1;  /* OR,C,A */
                {8'h61,8'h63} : dec_pc_inc2 = 1'b1;  /* OR,B,A */
                {8'h61,8'h64} : dec_pc_inc2 = 1'b1;  /* OR,E,A */
                {8'h61,8'h65} : dec_pc_inc2 = 1'b1;  /* OR,D,A */
                {8'h61,8'h66} : dec_pc_inc2 = 1'b1;  /* OR,L,A */
                {8'h61,8'h67} : dec_pc_inc2 = 1'b1;  /* OR,H,A */
                {8'h6b,8'hxx} : dec_pc_inc2 = 1'b1;  /* OR,A,saddr */
                {8'h6e,8'hxx} : dec_pc_inc2 = 1'b1;  /* OR,A,[HL+byte] */
                {8'h61,8'he0} : dec_pc_inc2 = 1'b1;  /* OR,A,[HL+B] */
                {8'h61,8'he2} : dec_pc_inc2 = 1'b1;  /* OR,A,[HL+C] */
                {8'h7c,8'hxx} : dec_pc_inc2 = 1'b1;  /* XOR,A,#byte */
                {8'h61,8'h78} : dec_pc_inc2 = 1'b1;  /* XOR,A,X */
                {8'h61,8'h7a} : dec_pc_inc2 = 1'b1;  /* XOR,A,C */
                {8'h61,8'h7b} : dec_pc_inc2 = 1'b1;  /* XOR,A,B */
                {8'h61,8'h7c} : dec_pc_inc2 = 1'b1;  /* XOR,A,E */
                {8'h61,8'h7d} : dec_pc_inc2 = 1'b1;  /* XOR,A,D */
                {8'h61,8'h7e} : dec_pc_inc2 = 1'b1;  /* XOR,A,L */
                {8'h61,8'h7f} : dec_pc_inc2 = 1'b1;  /* XOR,A,H */
                {8'h61,8'h70} : dec_pc_inc2 = 1'b1;  /* XOR,X,A */
                {8'h61,8'h71} : dec_pc_inc2 = 1'b1;  /* XOR,A,A */
                {8'h61,8'h72} : dec_pc_inc2 = 1'b1;  /* XOR,C,A */
                {8'h61,8'h73} : dec_pc_inc2 = 1'b1;  /* XOR,B,A */
                {8'h61,8'h74} : dec_pc_inc2 = 1'b1;  /* XOR,E,A */
                {8'h61,8'h75} : dec_pc_inc2 = 1'b1;  /* XOR,D,A */
                {8'h61,8'h76} : dec_pc_inc2 = 1'b1;  /* XOR,L,A */
                {8'h61,8'h77} : dec_pc_inc2 = 1'b1;  /* XOR,H,A */
                {8'h7b,8'hxx} : dec_pc_inc2 = 1'b1;  /* XOR,A,saddr */
                {8'h7e,8'hxx} : dec_pc_inc2 = 1'b1;  /* XOR,A,[HL+byte] */
                {8'h61,8'hf0} : dec_pc_inc2 = 1'b1;  /* XOR,A,[HL+B] */
                {8'h61,8'hf2} : dec_pc_inc2 = 1'b1;  /* XOR,A,[HL+C] */
                {8'h4c,8'hxx} : dec_pc_inc2 = 1'b1;  /* CMP,A,#byte */
                {8'h61,8'h48} : dec_pc_inc2 = 1'b1;  /* CMP,A,X */
                {8'h61,8'h4a} : dec_pc_inc2 = 1'b1;  /* CMP,A,C */
                {8'h61,8'h4b} : dec_pc_inc2 = 1'b1;  /* CMP,A,B */
                {8'h61,8'h4c} : dec_pc_inc2 = 1'b1;  /* CMP,A,E */
                {8'h61,8'h4d} : dec_pc_inc2 = 1'b1;  /* CMP,A,D */
                {8'h61,8'h4e} : dec_pc_inc2 = 1'b1;  /* CMP,A,L */
                {8'h61,8'h4f} : dec_pc_inc2 = 1'b1;  /* CMP,A,H */
                {8'h61,8'h40} : dec_pc_inc2 = 1'b1;  /* CMP,X,A */
                {8'h61,8'h41} : dec_pc_inc2 = 1'b1;  /* CMP,A,A */
                {8'h61,8'h42} : dec_pc_inc2 = 1'b1;  /* CMP,C,A */
                {8'h61,8'h43} : dec_pc_inc2 = 1'b1;  /* CMP,B,A */
                {8'h61,8'h44} : dec_pc_inc2 = 1'b1;  /* CMP,E,A */
                {8'h61,8'h45} : dec_pc_inc2 = 1'b1;  /* CMP,D,A */
                {8'h61,8'h46} : dec_pc_inc2 = 1'b1;  /* CMP,L,A */
                {8'h61,8'h47} : dec_pc_inc2 = 1'b1;  /* CMP,H,A */
                {8'h4b,8'hxx} : dec_pc_inc2 = 1'b1;  /* CMP,A,saddr */
                {8'h4e,8'hxx} : dec_pc_inc2 = 1'b1;  /* CMP,A,[HL+byte] */
                {8'h61,8'hc0} : dec_pc_inc2 = 1'b1;  /* CMP,A,[HL+B] */
                {8'h61,8'hc2} : dec_pc_inc2 = 1'b1;  /* CMP,A,[HL+C] */
                {8'hd4,8'hxx} : dec_pc_inc2 = 1'b1;  /* CMP0,,saddr */
                {8'h06,8'hxx} : dec_pc_inc2 = 1'b1;  /* ADDW,AX,saddrp */
                {8'h26,8'hxx} : dec_pc_inc2 = 1'b1;  /* SUBW,AX,saddrp */
                {8'h46,8'hxx} : dec_pc_inc2 = 1'b1;  /* CMPW,AX,saddrp */
                {8'ha4,8'hxx} : dec_pc_inc2 = 1'b1;  /* INC,,saddr */
                {8'hb4,8'hxx} : dec_pc_inc2 = 1'b1;  /* DEC,,saddr */
                {8'ha6,8'hxx} : dec_pc_inc2 = 1'b1;  /* INCW,,saddrp */
                {8'hb6,8'hxx} : dec_pc_inc2 = 1'b1;  /* DECW,,saddrp */
                {8'h31,8'h0a} : dec_pc_inc2 = 1'b1;  /* SHR,A,0 */
                {8'h31,8'h1a} : dec_pc_inc2 = 1'b1;  /* SHR,A,1 */
                {8'h31,8'h2a} : dec_pc_inc2 = 1'b1;  /* SHR,A,2 */
                {8'h31,8'h3a} : dec_pc_inc2 = 1'b1;  /* SHR,A,3 */
                {8'h31,8'h4a} : dec_pc_inc2 = 1'b1;  /* SHR,A,4 */
                {8'h31,8'h5a} : dec_pc_inc2 = 1'b1;  /* SHR,A,5 */
                {8'h31,8'h6a} : dec_pc_inc2 = 1'b1;  /* SHR,A,6 */
                {8'h31,8'h7a} : dec_pc_inc2 = 1'b1;  /* SHR,A,7 */
                {8'h31,8'h0e} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,0 */
                {8'h31,8'h1e} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,1 */
                {8'h31,8'h2e} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,2 */
                {8'h31,8'h3e} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,3 */
                {8'h31,8'h4e} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,4 */
                {8'h31,8'h5e} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,5 */
                {8'h31,8'h6e} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,6 */
                {8'h31,8'h7e} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,7 */
                {8'h31,8'h8e} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,8 */
                {8'h31,8'h9e} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,9 */
                {8'h31,8'hae} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,10 */
                {8'h31,8'hbe} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,11 */
                {8'h31,8'hce} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,12 */
                {8'h31,8'hde} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,13 */
                {8'h31,8'hee} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,14 */
                {8'h31,8'hfe} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,15 */
                {8'h31,8'h09} : dec_pc_inc2 = 1'b1;  /* SHL,A,0 */
                {8'h31,8'h19} : dec_pc_inc2 = 1'b1;  /* SHL,A,1 */
                {8'h31,8'h29} : dec_pc_inc2 = 1'b1;  /* SHL,A,2 */
                {8'h31,8'h39} : dec_pc_inc2 = 1'b1;  /* SHL,A,3 */
                {8'h31,8'h49} : dec_pc_inc2 = 1'b1;  /* SHL,A,4 */
                {8'h31,8'h59} : dec_pc_inc2 = 1'b1;  /* SHL,A,5 */
                {8'h31,8'h69} : dec_pc_inc2 = 1'b1;  /* SHL,A,6 */
                {8'h31,8'h79} : dec_pc_inc2 = 1'b1;  /* SHL,A,7 */
                {8'h31,8'h08} : dec_pc_inc2 = 1'b1;  /* SHL,B,0 */
                {8'h31,8'h18} : dec_pc_inc2 = 1'b1;  /* SHL,B,1 */
                {8'h31,8'h28} : dec_pc_inc2 = 1'b1;  /* SHL,B,2 */
                {8'h31,8'h38} : dec_pc_inc2 = 1'b1;  /* SHL,B,3 */
                {8'h31,8'h48} : dec_pc_inc2 = 1'b1;  /* SHL,B,4 */
                {8'h31,8'h58} : dec_pc_inc2 = 1'b1;  /* SHL,B,5 */
                {8'h31,8'h68} : dec_pc_inc2 = 1'b1;  /* SHL,B,6 */
                {8'h31,8'h78} : dec_pc_inc2 = 1'b1;  /* SHL,B,7 */
                {8'h31,8'h07} : dec_pc_inc2 = 1'b1;  /* SHL,C,0 */
                {8'h31,8'h17} : dec_pc_inc2 = 1'b1;  /* SHL,C,1 */
                {8'h31,8'h27} : dec_pc_inc2 = 1'b1;  /* SHL,C,2 */
                {8'h31,8'h37} : dec_pc_inc2 = 1'b1;  /* SHL,C,3 */
                {8'h31,8'h47} : dec_pc_inc2 = 1'b1;  /* SHL,C,4 */
                {8'h31,8'h57} : dec_pc_inc2 = 1'b1;  /* SHL,C,5 */
                {8'h31,8'h67} : dec_pc_inc2 = 1'b1;  /* SHL,C,6 */
                {8'h31,8'h77} : dec_pc_inc2 = 1'b1;  /* SHL,C,7 */
                {8'h31,8'h0d} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,0 */
                {8'h31,8'h1d} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,1 */
                {8'h31,8'h2d} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,2 */
                {8'h31,8'h3d} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,3 */
                {8'h31,8'h4d} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,4 */
                {8'h31,8'h5d} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,5 */
                {8'h31,8'h6d} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,6 */
                {8'h31,8'h7d} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,7 */
                {8'h31,8'h8d} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,8 */
                {8'h31,8'h9d} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,9 */
                {8'h31,8'had} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,10 */
                {8'h31,8'hbd} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,11 */
                {8'h31,8'hcd} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,12 */
                {8'h31,8'hdd} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,13 */
                {8'h31,8'hed} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,14 */
                {8'h31,8'hfd} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,15 */
                {8'h31,8'h0c} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,0 */
                {8'h31,8'h1c} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,1 */
                {8'h31,8'h2c} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,2 */
                {8'h31,8'h3c} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,3 */
                {8'h31,8'h4c} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,4 */
                {8'h31,8'h5c} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,5 */
                {8'h31,8'h6c} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,6 */
                {8'h31,8'h7c} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,7 */
                {8'h31,8'h8c} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,8 */
                {8'h31,8'h9c} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,9 */
                {8'h31,8'hac} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,10 */
                {8'h31,8'hbc} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,11 */
                {8'h31,8'hcc} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,12 */
                {8'h31,8'hdc} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,13 */
                {8'h31,8'hec} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,14 */
                {8'h31,8'hfc} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,15 */
                {8'h31,8'h0b} : dec_pc_inc2 = 1'b1;  /* SAR,A,0 */
                {8'h31,8'h1b} : dec_pc_inc2 = 1'b1;  /* SAR,A,1 */
                {8'h31,8'h2b} : dec_pc_inc2 = 1'b1;  /* SAR,A,2 */
                {8'h31,8'h3b} : dec_pc_inc2 = 1'b1;  /* SAR,A,3 */
                {8'h31,8'h4b} : dec_pc_inc2 = 1'b1;  /* SAR,A,4 */
                {8'h31,8'h5b} : dec_pc_inc2 = 1'b1;  /* SAR,A,5 */
                {8'h31,8'h6b} : dec_pc_inc2 = 1'b1;  /* SAR,A,6 */
                {8'h31,8'h7b} : dec_pc_inc2 = 1'b1;  /* SAR,A,7 */
                {8'h31,8'h0f} : dec_pc_inc2 = 1'b1;  /* SARW,AX,0 */
                {8'h31,8'h1f} : dec_pc_inc2 = 1'b1;  /* SARW,AX,1 */
                {8'h31,8'h2f} : dec_pc_inc2 = 1'b1;  /* SARW,AX,2 */
                {8'h31,8'h3f} : dec_pc_inc2 = 1'b1;  /* SARW,AX,3 */
                {8'h31,8'h4f} : dec_pc_inc2 = 1'b1;  /* SARW,AX,4 */
                {8'h31,8'h5f} : dec_pc_inc2 = 1'b1;  /* SARW,AX,5 */
                {8'h31,8'h6f} : dec_pc_inc2 = 1'b1;  /* SARW,AX,6 */
                {8'h31,8'h7f} : dec_pc_inc2 = 1'b1;  /* SARW,AX,7 */
                {8'h31,8'h8f} : dec_pc_inc2 = 1'b1;  /* SARW,AX,8 */
                {8'h31,8'h9f} : dec_pc_inc2 = 1'b1;  /* SARW,AX,9 */
                {8'h31,8'haf} : dec_pc_inc2 = 1'b1;  /* SARW,AX,10 */
                {8'h31,8'hbf} : dec_pc_inc2 = 1'b1;  /* SARW,AX,11 */
                {8'h31,8'hcf} : dec_pc_inc2 = 1'b1;  /* SARW,AX,12 */
                {8'h31,8'hdf} : dec_pc_inc2 = 1'b1;  /* SARW,AX,13 */
                {8'h31,8'hef} : dec_pc_inc2 = 1'b1;  /* SARW,AX,14 */
                {8'h31,8'hff} : dec_pc_inc2 = 1'b1;  /* SARW,AX,15 */
                {8'h61,8'hdb} : dec_pc_inc2 = 1'b1;  /* ROR,A,1 */
                {8'h61,8'heb} : dec_pc_inc2 = 1'b1;  /* ROL,A,1 */
                {8'h61,8'hfb} : dec_pc_inc2 = 1'b1;  /* RORC,A,1 */
                {8'h61,8'hdc} : dec_pc_inc2 = 1'b1;  /* ROLC,A,1 */
                {8'h61,8'hee} : dec_pc_inc2 = 1'b1;  /* ROLWC,AX,1 */
                {8'h61,8'hfe} : dec_pc_inc2 = 1'b1;  /* ROLWC,BC,1 */
                {8'h71,8'h8c} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,A.0 */
                {8'h71,8'h9c} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,A.1 */
                {8'h71,8'hac} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,A.2 */
                {8'h71,8'hbc} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,A.3 */
                {8'h71,8'hcc} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,A.4 */
                {8'h71,8'hdc} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,A.5 */
                {8'h71,8'hec} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,A.6 */
                {8'h71,8'hfc} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,A.7 */
                {8'h71,8'h84} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,[HL].0 */
                {8'h71,8'h94} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,[HL].1 */
                {8'h71,8'ha4} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,[HL].2 */
                {8'h71,8'hb4} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,[HL].3 */
                {8'h71,8'hc4} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,[HL].4 */
                {8'h71,8'hd4} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,[HL].5 */
                {8'h71,8'he4} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,[HL].6 */
                {8'h71,8'hf4} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,[HL].7 */
                {8'h71,8'h89} : dec_pc_inc2 = 1'b1;  /* MOV1,A.0,CY */
                {8'h71,8'h99} : dec_pc_inc2 = 1'b1;  /* MOV1,A.1,CY */
                {8'h71,8'ha9} : dec_pc_inc2 = 1'b1;  /* MOV1,A.2,CY */
                {8'h71,8'hb9} : dec_pc_inc2 = 1'b1;  /* MOV1,A.3,CY */
                {8'h71,8'hc9} : dec_pc_inc2 = 1'b1;  /* MOV1,A.4,CY */
                {8'h71,8'hd9} : dec_pc_inc2 = 1'b1;  /* MOV1,A.5,CY */
                {8'h71,8'he9} : dec_pc_inc2 = 1'b1;  /* MOV1,A.6,CY */
                {8'h71,8'hf9} : dec_pc_inc2 = 1'b1;  /* MOV1,A.7,CY */
                {8'h71,8'h81} : dec_pc_inc2 = 1'b1;  /* MOV1,[HL].0,CY */
                {8'h71,8'h91} : dec_pc_inc2 = 1'b1;  /* MOV1,[HL].1,CY */
                {8'h71,8'ha1} : dec_pc_inc2 = 1'b1;  /* MOV1,[HL].2,CY */
                {8'h71,8'hb1} : dec_pc_inc2 = 1'b1;  /* MOV1,[HL].3,CY */
                {8'h71,8'hc1} : dec_pc_inc2 = 1'b1;  /* MOV1,[HL].4,CY */
                {8'h71,8'hd1} : dec_pc_inc2 = 1'b1;  /* MOV1,[HL].5,CY */
                {8'h71,8'he1} : dec_pc_inc2 = 1'b1;  /* MOV1,[HL].6,CY */
                {8'h71,8'hf1} : dec_pc_inc2 = 1'b1;  /* MOV1,[HL].7,CY */
                {8'h71,8'h8d} : dec_pc_inc2 = 1'b1;  /* AND1,CY,A.0 */
                {8'h71,8'h9d} : dec_pc_inc2 = 1'b1;  /* AND1,CY,A.1 */
                {8'h71,8'had} : dec_pc_inc2 = 1'b1;  /* AND1,CY,A.2 */
                {8'h71,8'hbd} : dec_pc_inc2 = 1'b1;  /* AND1,CY,A.3 */
                {8'h71,8'hcd} : dec_pc_inc2 = 1'b1;  /* AND1,CY,A.4 */
                {8'h71,8'hdd} : dec_pc_inc2 = 1'b1;  /* AND1,CY,A.5 */
                {8'h71,8'hed} : dec_pc_inc2 = 1'b1;  /* AND1,CY,A.6 */
                {8'h71,8'hfd} : dec_pc_inc2 = 1'b1;  /* AND1,CY,A.7 */
                {8'h71,8'h85} : dec_pc_inc2 = 1'b1;  /* AND1,CY,[HL].0 */
                {8'h71,8'h95} : dec_pc_inc2 = 1'b1;  /* AND1,CY,[HL].1 */
                {8'h71,8'ha5} : dec_pc_inc2 = 1'b1;  /* AND1,CY,[HL].2 */
                {8'h71,8'hb5} : dec_pc_inc2 = 1'b1;  /* AND1,CY,[HL].3 */
                {8'h71,8'hc5} : dec_pc_inc2 = 1'b1;  /* AND1,CY,[HL].4 */
                {8'h71,8'hd5} : dec_pc_inc2 = 1'b1;  /* AND1,CY,[HL].5 */
                {8'h71,8'he5} : dec_pc_inc2 = 1'b1;  /* AND1,CY,[HL].6 */
                {8'h71,8'hf5} : dec_pc_inc2 = 1'b1;  /* AND1,CY,[HL].7 */
                {8'h71,8'h8e} : dec_pc_inc2 = 1'b1;  /* OR1,CY,A.0 */
                {8'h71,8'h9e} : dec_pc_inc2 = 1'b1;  /* OR1,CY,A.1 */
                {8'h71,8'hae} : dec_pc_inc2 = 1'b1;  /* OR1,CY,A.2 */
                {8'h71,8'hbe} : dec_pc_inc2 = 1'b1;  /* OR1,CY,A.3 */
                {8'h71,8'hce} : dec_pc_inc2 = 1'b1;  /* OR1,CY,A.4 */
                {8'h71,8'hde} : dec_pc_inc2 = 1'b1;  /* OR1,CY,A.5 */
                {8'h71,8'hee} : dec_pc_inc2 = 1'b1;  /* OR1,CY,A.6 */
                {8'h71,8'hfe} : dec_pc_inc2 = 1'b1;  /* OR1,CY,A.7 */
                {8'h71,8'h86} : dec_pc_inc2 = 1'b1;  /* OR1,CY,[HL].0 */
                {8'h71,8'h96} : dec_pc_inc2 = 1'b1;  /* OR1,CY,[HL].1 */
                {8'h71,8'ha6} : dec_pc_inc2 = 1'b1;  /* OR1,CY,[HL].2 */
                {8'h71,8'hb6} : dec_pc_inc2 = 1'b1;  /* OR1,CY,[HL].3 */
                {8'h71,8'hc6} : dec_pc_inc2 = 1'b1;  /* OR1,CY,[HL].4 */
                {8'h71,8'hd6} : dec_pc_inc2 = 1'b1;  /* OR1,CY,[HL].5 */
                {8'h71,8'he6} : dec_pc_inc2 = 1'b1;  /* OR1,CY,[HL].6 */
                {8'h71,8'hf6} : dec_pc_inc2 = 1'b1;  /* OR1,CY,[HL].7 */
                {8'h71,8'h8f} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,A.0 */
                {8'h71,8'h9f} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,A.1 */
                {8'h71,8'haf} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,A.2 */
                {8'h71,8'hbf} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,A.3 */
                {8'h71,8'hcf} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,A.4 */
                {8'h71,8'hdf} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,A.5 */
                {8'h71,8'hef} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,A.6 */
                {8'h71,8'hff} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,A.7 */
                {8'h71,8'h87} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,[HL].0 */
                {8'h71,8'h97} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,[HL].1 */
                {8'h71,8'ha7} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,[HL].2 */
                {8'h71,8'hb7} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,[HL].3 */
                {8'h71,8'hc7} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,[HL].4 */
                {8'h71,8'hd7} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,[HL].5 */
                {8'h71,8'he7} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,[HL].6 */
                {8'h71,8'hf7} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,[HL].7 */
                {8'h71,8'h8a} : dec_pc_inc2 = 1'b1;  /* SET1,,A.0 */
                {8'h71,8'h9a} : dec_pc_inc2 = 1'b1;  /* SET1,,A.1 */
                {8'h71,8'haa} : dec_pc_inc2 = 1'b1;  /* SET1,,A.2 */
                {8'h71,8'hba} : dec_pc_inc2 = 1'b1;  /* SET1,,A.3 */
                {8'h71,8'hca} : dec_pc_inc2 = 1'b1;  /* SET1,,A.4 */
                {8'h71,8'hda} : dec_pc_inc2 = 1'b1;  /* SET1,,A.5 */
                {8'h71,8'hea} : dec_pc_inc2 = 1'b1;  /* SET1,,A.6 */
                {8'h71,8'hfa} : dec_pc_inc2 = 1'b1;  /* SET1,,A.7 */
                {8'h71,8'h82} : dec_pc_inc2 = 1'b1;  /* SET1,,[HL].0 */
                {8'h71,8'h92} : dec_pc_inc2 = 1'b1;  /* SET1,,[HL].1 */
                {8'h71,8'ha2} : dec_pc_inc2 = 1'b1;  /* SET1,,[HL].2 */
                {8'h71,8'hb2} : dec_pc_inc2 = 1'b1;  /* SET1,,[HL].3 */
                {8'h71,8'hc2} : dec_pc_inc2 = 1'b1;  /* SET1,,[HL].4 */
                {8'h71,8'hd2} : dec_pc_inc2 = 1'b1;  /* SET1,,[HL].5 */
                {8'h71,8'he2} : dec_pc_inc2 = 1'b1;  /* SET1,,[HL].6 */
                {8'h71,8'hf2} : dec_pc_inc2 = 1'b1;  /* SET1,,[HL].7 */
                {8'h71,8'h8b} : dec_pc_inc2 = 1'b1;  /* CLR1,,A.0 */
                {8'h71,8'h9b} : dec_pc_inc2 = 1'b1;  /* CLR1,,A.1 */
                {8'h71,8'hab} : dec_pc_inc2 = 1'b1;  /* CLR1,,A.2 */
                {8'h71,8'hbb} : dec_pc_inc2 = 1'b1;  /* CLR1,,A.3 */
                {8'h71,8'hcb} : dec_pc_inc2 = 1'b1;  /* CLR1,,A.4 */
                {8'h71,8'hdb} : dec_pc_inc2 = 1'b1;  /* CLR1,,A.5 */
                {8'h71,8'heb} : dec_pc_inc2 = 1'b1;  /* CLR1,,A.6 */
                {8'h71,8'hfb} : dec_pc_inc2 = 1'b1;  /* CLR1,,A.7 */
                {8'h71,8'h83} : dec_pc_inc2 = 1'b1;  /* CLR1,,[HL].0 */
                {8'h71,8'h93} : dec_pc_inc2 = 1'b1;  /* CLR1,,[HL].1 */
                {8'h71,8'ha3} : dec_pc_inc2 = 1'b1;  /* CLR1,,[HL].2 */
                {8'h71,8'hb3} : dec_pc_inc2 = 1'b1;  /* CLR1,,[HL].3 */
                {8'h71,8'hc3} : dec_pc_inc2 = 1'b1;  /* CLR1,,[HL].4 */
                {8'h71,8'hd3} : dec_pc_inc2 = 1'b1;  /* CLR1,,[HL].5 */
                {8'h71,8'he3} : dec_pc_inc2 = 1'b1;  /* CLR1,,[HL].6 */
                {8'h71,8'hf3} : dec_pc_inc2 = 1'b1;  /* CLR1,,[HL].7 */
                {8'h71,8'h80} : dec_pc_inc2 = 1'b1;  /* SET1,,CY */
                {8'h71,8'h88} : dec_pc_inc2 = 1'b1;  /* CLR1,,CY */
                {8'h71,8'hc0} : dec_pc_inc2 = 1'b1;  /* NOT1,,CY */
                {8'h61,8'hca} : dec_pc_inc2 = 1'b1;  /* CALL,,AX */
                {8'h61,8'hda} : dec_pc_inc2 = 1'b1;  /* CALL,,BC */
                {8'h61,8'hea} : dec_pc_inc2 = 1'b1;  /* CALL,,DE */
                {8'h61,8'hfa} : dec_pc_inc2 = 1'b1;  /* CALL,,HL */
                {8'h61,8'h84} : dec_pc_inc2 = 1'b1;  /* CALLT,,[0080h] */
                {8'h61,8'h94} : dec_pc_inc2 = 1'b1;  /* CALLT,,[0082h] */
                {8'h61,8'ha4} : dec_pc_inc2 = 1'b1;  /* CALLT,,[0084h] */
                {8'h61,8'hb4} : dec_pc_inc2 = 1'b1;  /* CALLT,,[0086h] */
                {8'h61,8'hc4} : dec_pc_inc2 = 1'b1;  /* CALLT,,[0088h] */
                {8'h61,8'hd4} : dec_pc_inc2 = 1'b1;  /* CALLT,,[008Ah] */
                {8'h61,8'he4} : dec_pc_inc2 = 1'b1;  /* CALLT,,[008Ch] */
                {8'h61,8'hf4} : dec_pc_inc2 = 1'b1;  /* CALLT,,[008Eh] */
                {8'h61,8'h85} : dec_pc_inc2 = 1'b1;  /* CALLT,,[0090h] */
                {8'h61,8'h95} : dec_pc_inc2 = 1'b1;  /* CALLT,,[0092h] */
                {8'h61,8'ha5} : dec_pc_inc2 = 1'b1;  /* CALLT,,[0094h] */
                {8'h61,8'hb5} : dec_pc_inc2 = 1'b1;  /* CALLT,,[0096h] */
                {8'h61,8'hc5} : dec_pc_inc2 = 1'b1;  /* CALLT,,[0098h] */
                {8'h61,8'hd5} : dec_pc_inc2 = 1'b1;  /* CALLT,,[009Ah] */
                {8'h61,8'he5} : dec_pc_inc2 = 1'b1;  /* CALLT,,[009Ch] */
                {8'h61,8'hf5} : dec_pc_inc2 = 1'b1;  /* CALLT,,[009Eh] */
                {8'h61,8'h86} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00A0h] */
                {8'h61,8'h96} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00A2h] */
                {8'h61,8'ha6} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00A4h] */
                {8'h61,8'hb6} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00A6h] */
                {8'h61,8'hc6} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00A8h] */
                {8'h61,8'hd6} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00AAh] */
                {8'h61,8'he6} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00ACh] */
                {8'h61,8'hf6} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00AEh] */
                {8'h61,8'h87} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00B0h] */
                {8'h61,8'h97} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00B2h] */
                {8'h61,8'ha7} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00B4h] */
                {8'h61,8'hb7} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00B6h] */
                {8'h61,8'hc7} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00B8h] */
                {8'h61,8'hd7} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00BAh] */
                {8'h61,8'he7} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00BCh] */
                {8'h61,8'hf7} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00BEh] */
                {8'h61,8'hcc} : dec_pc_inc2 = 1'b1;  /* BRK,, */
                {8'h61,8'hec} : dec_pc_inc2 = 1'b1;  /* RETB,, */
                {8'h61,8'hfc} : dec_pc_inc2 = 1'b1;  /* RETI,, */
                {8'h61,8'hdd} : dec_pc_inc2 = 1'b1;  /* PUSH,,PSW */
                {8'h61,8'hcd} : dec_pc_inc2 = 1'b1;  /* POP,,PSW */
                {8'h10,8'hxx} : dec_pc_inc2 = 1'b1;  /* ADDW,SP,#byte */
                {8'h20,8'hxx} : dec_pc_inc2 = 1'b1;  /* SUBW,SP,#byte */
                {8'hef,8'hxx} : dec_pc_inc2 = 1'b1;  /* BR,,$addr8 */
                {8'h61,8'hcb} : dec_pc_inc2 = 1'b1;  /* BR,,AX */
                {8'hdc,8'hxx} : dec_pc_inc2 = 1'b1;  /* BC,,$addr8 */
                {8'hde,8'hxx} : dec_pc_inc2 = 1'b1;  /* BNC,,$addr8 */
                {8'hdd,8'hxx} : dec_pc_inc2 = 1'b1;  /* BZ,,$addr8 */
                {8'hdf,8'hxx} : dec_pc_inc2 = 1'b1;  /* BNZ,,$addr8 */
                {8'h61,8'hc8} : dec_pc_inc2 = 1'b1;  /* SKC,, */
                {8'h61,8'hd8} : dec_pc_inc2 = 1'b1;  /* SKNC,, */
                {8'h61,8'he8} : dec_pc_inc2 = 1'b1;  /* SKZ,, */
                {8'h61,8'hf8} : dec_pc_inc2 = 1'b1;  /* SKNZ,, */
                {8'h61,8'he3} : dec_pc_inc2 = 1'b1;  /* SKH,, */
                {8'h61,8'hf3} : dec_pc_inc2 = 1'b1;  /* SKNH,, */
                {8'h61,8'hcf} : dec_pc_inc2 = 1'b1;  /* SEL,,RB0 */
                {8'h61,8'hdf} : dec_pc_inc2 = 1'b1;  /* SEL,,RB1 */
                {8'h61,8'hef} : dec_pc_inc2 = 1'b1;  /* SEL,,RB2 */
                {8'h61,8'hff} : dec_pc_inc2 = 1'b1;  /* SEL,,RB3 */
                {8'h61,8'hed} : dec_pc_inc2 = 1'b1;  /* HALT,, */
                {8'h61,8'hfd} : dec_pc_inc2 = 1'b1;  /* STOP,, */
                {8'h61,8'ha1} : dec_pc_inc2 = 1'b1;  /* SOFT2,,BREAK */
                {8'h61,8'h81} : dec_pc_inc2 = 1'b1;  /* ALT1,, */
                {8'h61,8'h91} : dec_pc_inc2 = 1'b1;  /* ALT2,, */
                {8'h61,8'h88} : dec_pc_inc2 = 1'b1;  /* XCH,A,X */
                {8'h61,8'h98} : dec_pc_inc2 = 1'b1;  /* XCH,A,X */
                {8'h61,8'h99} : dec_pc_inc2 = 1'b1;  /* XCH,A,X */
                {8'h61,8'h9a} : dec_pc_inc2 = 1'b1;  /* XCH,A,C */
                {8'h61,8'h9b} : dec_pc_inc2 = 1'b1;  /* XCH,A,B */
                {8'h61,8'h9c} : dec_pc_inc2 = 1'b1;  /* XCH,A,E */
                {8'h61,8'h9d} : dec_pc_inc2 = 1'b1;  /* XCH,A,D */
                {8'h61,8'h9e} : dec_pc_inc2 = 1'b1;  /* XCH,A,L */
                {8'h61,8'h9f} : dec_pc_inc2 = 1'b1;  /* XCH,A,H */
                {8'h61,8'hbe} : dec_pc_inc2 = 1'b1;  /* XCH,A,[DE] */
                {8'h61,8'hbc} : dec_pc_inc2 = 1'b1;  /* XCH,A,[HL] */
                {8'h61,8'h19} : dec_pc_inc2 = 1'b1;  /* ADDC,A,A */
                {8'h61,8'h39} : dec_pc_inc2 = 1'b1;  /* SUBC,A,A */
                {8'h61,8'hd1} : dec_pc_inc2 = 1'b1;  /* AND,A,[HL+B] */
                {8'h61,8'he1} : dec_pc_inc2 = 1'b1;  /* OR,A,[HL+B] */
                {8'h61,8'hf1} : dec_pc_inc2 = 1'b1;  /* XOR,A,[HL+B] */
                {8'h61,8'h83} : dec_pc_inc2 = 1'b1;  /* ADD,A,[HL+C] */
                {8'h61,8'h93} : dec_pc_inc2 = 1'b1;  /* ADDC,A,[HL+C] */
                {8'h61,8'ha3} : dec_pc_inc2 = 1'b1;  /* SUB,A,[HL+C] */
                {8'h61,8'hb3} : dec_pc_inc2 = 1'b1;  /* SUBC,A,[HL+C] */
                {8'h71,8'h90} : dec_pc_inc2 = 1'b1;  /* SET1,,CY */
                {8'h71,8'ha0} : dec_pc_inc2 = 1'b1;  /* SET1,,CY */
                {8'h71,8'hb0} : dec_pc_inc2 = 1'b1;  /* SET1,,CY */
                {8'h71,8'hd0} : dec_pc_inc2 = 1'b1;  /* NOT1,,CY */
                {8'h71,8'he0} : dec_pc_inc2 = 1'b1;  /* NOT1,,CY */
                {8'h71,8'hf0} : dec_pc_inc2 = 1'b1;  /* NOT1,,CY */
                {8'h71,8'h98} : dec_pc_inc2 = 1'b1;  /* CLR1,,CY */
                {8'h71,8'ha8} : dec_pc_inc2 = 1'b1;  /* CLR1,,CY */
                {8'h71,8'hb8} : dec_pc_inc2 = 1'b1;  /* CLR1,,CY */
                {8'h71,8'hc8} : dec_pc_inc2 = 1'b1;  /* NOT1,,CY */
                {8'h71,8'hd8} : dec_pc_inc2 = 1'b1;  /* NOT1,,CY */
                {8'h71,8'he8} : dec_pc_inc2 = 1'b1;  /* NOT1,,CY */
                {8'h71,8'hf8} : dec_pc_inc2 = 1'b1;  /* NOT1,,CY */
                {8'h31,8'h8a} : dec_pc_inc2 = 1'b1;  /* SHR,A,0 */
                {8'h31,8'h9a} : dec_pc_inc2 = 1'b1;  /* SHR,A,1 */
                {8'h31,8'haa} : dec_pc_inc2 = 1'b1;  /* SHR,A,2 */
                {8'h31,8'hba} : dec_pc_inc2 = 1'b1;  /* SHR,A,3 */
                {8'h31,8'hca} : dec_pc_inc2 = 1'b1;  /* SHR,A,4 */
                {8'h31,8'hda} : dec_pc_inc2 = 1'b1;  /* SHR,A,5 */
                {8'h31,8'hea} : dec_pc_inc2 = 1'b1;  /* SHR,A,6 */
                {8'h31,8'hfa} : dec_pc_inc2 = 1'b1;  /* SHR,A,7 */
                {8'h31,8'h89} : dec_pc_inc2 = 1'b1;  /* SHL,A,0 */
                {8'h31,8'h99} : dec_pc_inc2 = 1'b1;  /* SHL,A,1 */
                {8'h31,8'ha9} : dec_pc_inc2 = 1'b1;  /* SHL,A,2 */
                {8'h31,8'hb9} : dec_pc_inc2 = 1'b1;  /* SHL,A,3 */
                {8'h31,8'hc9} : dec_pc_inc2 = 1'b1;  /* SHL,A,4 */
                {8'h31,8'hd9} : dec_pc_inc2 = 1'b1;  /* SHL,A,5 */
                {8'h31,8'he9} : dec_pc_inc2 = 1'b1;  /* SHL,A,6 */
                {8'h31,8'hf9} : dec_pc_inc2 = 1'b1;  /* SHL,A,7 */
                {8'h31,8'h88} : dec_pc_inc2 = 1'b1;  /* SHL,B,0 */
                {8'h31,8'h98} : dec_pc_inc2 = 1'b1;  /* SHL,B,1 */
                {8'h31,8'ha8} : dec_pc_inc2 = 1'b1;  /* SHL,B,2 */
                {8'h31,8'hb8} : dec_pc_inc2 = 1'b1;  /* SHL,B,3 */
                {8'h31,8'hc8} : dec_pc_inc2 = 1'b1;  /* SHL,B,4 */
                {8'h31,8'hd8} : dec_pc_inc2 = 1'b1;  /* SHL,B,5 */
                {8'h31,8'he8} : dec_pc_inc2 = 1'b1;  /* SHL,B,6 */
                {8'h31,8'hf8} : dec_pc_inc2 = 1'b1;  /* SHL,B,7 */
                {8'h31,8'h87} : dec_pc_inc2 = 1'b1;  /* SHL,C,0 */
                {8'h31,8'h97} : dec_pc_inc2 = 1'b1;  /* SHL,C,1 */
                {8'h31,8'ha7} : dec_pc_inc2 = 1'b1;  /* SHL,C,2 */
                {8'h31,8'hb7} : dec_pc_inc2 = 1'b1;  /* SHL,C,3 */
                {8'h31,8'hc7} : dec_pc_inc2 = 1'b1;  /* SHL,C,4 */
                {8'h31,8'hd7} : dec_pc_inc2 = 1'b1;  /* SHL,C,5 */
                {8'h31,8'he7} : dec_pc_inc2 = 1'b1;  /* SHL,C,6 */
                {8'h31,8'hf7} : dec_pc_inc2 = 1'b1;  /* SHL,C,7 */
                {8'h31,8'h8b} : dec_pc_inc2 = 1'b1;  /* SAR,A,0 */
                {8'h31,8'h9b} : dec_pc_inc2 = 1'b1;  /* SAR,A,1 */
                {8'h31,8'hab} : dec_pc_inc2 = 1'b1;  /* SAR,A,2 */
                {8'h31,8'hbb} : dec_pc_inc2 = 1'b1;  /* SAR,A,3 */
                {8'h31,8'hcb} : dec_pc_inc2 = 1'b1;  /* SAR,A,4 */
                {8'h31,8'hdb} : dec_pc_inc2 = 1'b1;  /* SAR,A,5 */
                {8'h31,8'heb} : dec_pc_inc2 = 1'b1;  /* SAR,A,6 */
                {8'h31,8'hfb} : dec_pc_inc2 = 1'b1;  /* SAR,A,7 */
                {8'h31,8'h06} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'h16} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'h26} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'h36} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'h46} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'h56} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'h66} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'h76} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'h86} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'h96} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'ha6} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'hb6} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'hc6} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'hd6} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'he6} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'hf6} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                default : dec_pc_inc2 = 1'b0;
            endcase
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h50,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,X,#byte */
                {8'h51,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,A,#byte */
                {8'h52,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,C,#byte */
                {8'h53,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,B,#byte */
                {8'h54,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,E,#byte */
                {8'h55,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,D,#byte */
                {8'h56,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,L,#byte */
                {8'h57,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,H,#byte */
                {8'h8d,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,A,saddr */
                {8'h9d,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,saddr,A */
                {8'h8e,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,A,sfr */
                {8'h9e,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,sfr,A */
                {8'h41,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,ES,#byte */
                {8'h8a,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,A,[DE+byte] */
                {8'h9a,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,[DE+byte],A */
                {8'h8c,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,A,[HL+byte] */
                {8'h9c,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,[HL+byte],A */
                {8'h61,8'hc9,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,A,[HL+B] */
                {8'h61,8'hd9,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,[HL+B],A */
                {8'h61,8'he9,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,A,[HL+C] */
                {8'h61,8'hf9,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,[HL+C],A */
                {8'h88,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,A,[SP+byte] */
                {8'h98,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,[SP+byte],A */
                {8'he8,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,B,saddr */
                {8'hf8,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,C,saddr */
                {8'hd8,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV,X,saddr */
                {8'h61,8'h8a,2'bxx} : dec_pc_inc2 = 1'b1;  /* XCH,A,C */
                {8'h61,8'h8b,2'bxx} : dec_pc_inc2 = 1'b1;  /* XCH,A,B */
                {8'h61,8'h8c,2'bxx} : dec_pc_inc2 = 1'b1;  /* XCH,A,E */
                {8'h61,8'h8d,2'bxx} : dec_pc_inc2 = 1'b1;  /* XCH,A,D */
                {8'h61,8'h8e,2'bxx} : dec_pc_inc2 = 1'b1;  /* XCH,A,L */
                {8'h61,8'h8f,2'bxx} : dec_pc_inc2 = 1'b1;  /* XCH,A,H */
                {8'h61,8'hae,2'bx1} : dec_pc_inc2 = 1'b1;  /* XCH,A,[DE] */
                {8'h61,8'hac,2'bx1} : dec_pc_inc2 = 1'b1;  /* XCH,A,[HL] */
                {8'h61,8'hb9,2'bx1} : dec_pc_inc2 = 1'b1;  /* XCH,A,[HL+B] */
                {8'h61,8'ha9,2'bx1} : dec_pc_inc2 = 1'b1;  /* XCH,A,[HL+C] */
                {8'he4,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* ONEB,,saddr */
                {8'hf4,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* CLRB,,saddr */
                {8'had,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOVW,AX,saddrp */
                {8'hbd,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOVW,saddrp,AX */
                {8'hae,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOVW,AX,sfrp */
                {8'hbe,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOVW,sfrp,AX */
                {8'haa,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOVW,AX,[DE+byte] */
                {8'hba,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOVW,[DE+byte],AX */
                {8'hac,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOVW,AX,[HL+byte] */
                {8'hbc,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOVW,[HL+byte],AX */
                {8'ha8,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOVW,AX,[SP+byte] */
                {8'hb8,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOVW,[SP+byte],AX */
                {8'hda,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOVW,BC,saddrp */
                {8'hea,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOVW,DE,saddrp */
                {8'hfa,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOVW,HL,saddrp */
                {8'h0c,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADD,A,#byte */
                {8'h61,8'h08,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADD,A,X */
                {8'h61,8'h0a,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADD,A,C */
                {8'h61,8'h0b,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADD,A,B */
                {8'h61,8'h0c,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADD,A,E */
                {8'h61,8'h0d,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADD,A,D */
                {8'h61,8'h0e,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADD,A,L */
                {8'h61,8'h0f,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADD,A,H */
                {8'h61,8'h00,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADD,X,A */
                {8'h61,8'h01,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADD,A,A */
                {8'h61,8'h02,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADD,C,A */
                {8'h61,8'h03,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADD,B,A */
                {8'h61,8'h04,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADD,E,A */
                {8'h61,8'h05,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADD,D,A */
                {8'h61,8'h06,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADD,L,A */
                {8'h61,8'h07,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADD,H,A */
                {8'h0b,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADD,A,saddr */
                {8'h0e,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADD,A,[HL+byte] */
                {8'h61,8'h80,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADD,A,[HL+B] */
                {8'h61,8'h82,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADD,A,[HL+C] */
                {8'h1c,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDC,A,#byte */
                {8'h61,8'h18,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDC,A,X */
                {8'h61,8'h1a,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDC,A,C */
                {8'h61,8'h1b,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDC,A,B */
                {8'h61,8'h1c,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDC,A,E */
                {8'h61,8'h1d,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDC,A,D */
                {8'h61,8'h1e,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDC,A,L */
                {8'h61,8'h1f,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDC,A,H */
                {8'h61,8'h10,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDC,X,A */
                {8'h61,8'h11,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDC,A,A */
                {8'h61,8'h12,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDC,C,A */
                {8'h61,8'h13,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDC,B,A */
                {8'h61,8'h14,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDC,E,A */
                {8'h61,8'h15,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDC,D,A */
                {8'h61,8'h16,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDC,L,A */
                {8'h61,8'h17,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDC,H,A */
                {8'h1b,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDC,A,saddr */
                {8'h1e,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDC,A,[HL+byte] */
                {8'h61,8'h90,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDC,A,[HL+B] */
                {8'h61,8'h92,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDC,A,[HL+C] */
                {8'h2c,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUB,A,#byte */
                {8'h61,8'h28,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUB,A,X */
                {8'h61,8'h2a,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUB,A,C */
                {8'h61,8'h2b,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUB,A,B */
                {8'h61,8'h2c,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUB,A,E */
                {8'h61,8'h2d,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUB,A,D */
                {8'h61,8'h2e,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUB,A,L */
                {8'h61,8'h2f,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUB,A,H */
                {8'h61,8'h20,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUB,X,A */
                {8'h61,8'h21,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUB,A,A */
                {8'h61,8'h22,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUB,C,A */
                {8'h61,8'h23,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUB,B,A */
                {8'h61,8'h24,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUB,E,A */
                {8'h61,8'h25,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUB,D,A */
                {8'h61,8'h26,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUB,L,A */
                {8'h61,8'h27,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUB,H,A */
                {8'h2b,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUB,A,saddr */
                {8'h2e,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUB,A,[HL+byte] */
                {8'h61,8'ha0,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUB,A,[HL+B] */
                {8'h61,8'ha2,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUB,A,[HL+C] */
                {8'h3c,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBC,A,#byte */
                {8'h61,8'h38,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBC,A,X */
                {8'h61,8'h3a,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBC,A,C */
                {8'h61,8'h3b,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBC,A,B */
                {8'h61,8'h3c,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBC,A,E */
                {8'h61,8'h3d,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBC,A,D */
                {8'h61,8'h3e,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBC,A,L */
                {8'h61,8'h3f,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBC,A,H */
                {8'h61,8'h30,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBC,X,A */
                {8'h61,8'h31,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBC,A,A */
                {8'h61,8'h32,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBC,C,A */
                {8'h61,8'h33,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBC,B,A */
                {8'h61,8'h34,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBC,E,A */
                {8'h61,8'h35,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBC,D,A */
                {8'h61,8'h36,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBC,L,A */
                {8'h61,8'h37,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBC,H,A */
                {8'h3b,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBC,A,saddr */
                {8'h3e,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBC,A,[HL+byte] */
                {8'h61,8'hb0,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBC,A,[HL+B] */
                {8'h61,8'hb2,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBC,A,[HL+C] */
                {8'h5c,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND,A,#byte */
                {8'h61,8'h58,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND,A,X */
                {8'h61,8'h5a,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND,A,C */
                {8'h61,8'h5b,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND,A,B */
                {8'h61,8'h5c,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND,A,E */
                {8'h61,8'h5d,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND,A,D */
                {8'h61,8'h5e,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND,A,L */
                {8'h61,8'h5f,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND,A,H */
                {8'h61,8'h50,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND,X,A */
                {8'h61,8'h51,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND,A,A */
                {8'h61,8'h52,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND,C,A */
                {8'h61,8'h53,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND,B,A */
                {8'h61,8'h54,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND,E,A */
                {8'h61,8'h55,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND,D,A */
                {8'h61,8'h56,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND,L,A */
                {8'h61,8'h57,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND,H,A */
                {8'h5b,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND,A,saddr */
                {8'h5e,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND,A,[HL+byte] */
                {8'h61,8'hd0,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND,A,[HL+B] */
                {8'h61,8'hd2,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND,A,[HL+C] */
                {8'h6c,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR,A,#byte */
                {8'h61,8'h68,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR,A,X */
                {8'h61,8'h6a,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR,A,C */
                {8'h61,8'h6b,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR,A,B */
                {8'h61,8'h6c,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR,A,E */
                {8'h61,8'h6d,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR,A,D */
                {8'h61,8'h6e,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR,A,L */
                {8'h61,8'h6f,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR,A,H */
                {8'h61,8'h60,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR,X,A */
                {8'h61,8'h61,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR,A,A */
                {8'h61,8'h62,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR,C,A */
                {8'h61,8'h63,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR,B,A */
                {8'h61,8'h64,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR,E,A */
                {8'h61,8'h65,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR,D,A */
                {8'h61,8'h66,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR,L,A */
                {8'h61,8'h67,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR,H,A */
                {8'h6b,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR,A,saddr */
                {8'h6e,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR,A,[HL+byte] */
                {8'h61,8'he0,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR,A,[HL+B] */
                {8'h61,8'he2,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR,A,[HL+C] */
                {8'h7c,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR,A,#byte */
                {8'h61,8'h78,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR,A,X */
                {8'h61,8'h7a,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR,A,C */
                {8'h61,8'h7b,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR,A,B */
                {8'h61,8'h7c,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR,A,E */
                {8'h61,8'h7d,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR,A,D */
                {8'h61,8'h7e,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR,A,L */
                {8'h61,8'h7f,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR,A,H */
                {8'h61,8'h70,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR,X,A */
                {8'h61,8'h71,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR,A,A */
                {8'h61,8'h72,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR,C,A */
                {8'h61,8'h73,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR,B,A */
                {8'h61,8'h74,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR,E,A */
                {8'h61,8'h75,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR,D,A */
                {8'h61,8'h76,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR,L,A */
                {8'h61,8'h77,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR,H,A */
                {8'h7b,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR,A,saddr */
                {8'h7e,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR,A,[HL+byte] */
                {8'h61,8'hf0,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR,A,[HL+B] */
                {8'h61,8'hf2,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR,A,[HL+C] */
                {8'h4c,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* CMP,A,#byte */
                {8'h61,8'h48,2'bxx} : dec_pc_inc2 = 1'b1;  /* CMP,A,X */
                {8'h61,8'h4a,2'bxx} : dec_pc_inc2 = 1'b1;  /* CMP,A,C */
                {8'h61,8'h4b,2'bxx} : dec_pc_inc2 = 1'b1;  /* CMP,A,B */
                {8'h61,8'h4c,2'bxx} : dec_pc_inc2 = 1'b1;  /* CMP,A,E */
                {8'h61,8'h4d,2'bxx} : dec_pc_inc2 = 1'b1;  /* CMP,A,D */
                {8'h61,8'h4e,2'bxx} : dec_pc_inc2 = 1'b1;  /* CMP,A,L */
                {8'h61,8'h4f,2'bxx} : dec_pc_inc2 = 1'b1;  /* CMP,A,H */
                {8'h61,8'h40,2'bxx} : dec_pc_inc2 = 1'b1;  /* CMP,X,A */
                {8'h61,8'h41,2'bxx} : dec_pc_inc2 = 1'b1;  /* CMP,A,A */
                {8'h61,8'h42,2'bxx} : dec_pc_inc2 = 1'b1;  /* CMP,C,A */
                {8'h61,8'h43,2'bxx} : dec_pc_inc2 = 1'b1;  /* CMP,B,A */
                {8'h61,8'h44,2'bxx} : dec_pc_inc2 = 1'b1;  /* CMP,E,A */
                {8'h61,8'h45,2'bxx} : dec_pc_inc2 = 1'b1;  /* CMP,D,A */
                {8'h61,8'h46,2'bxx} : dec_pc_inc2 = 1'b1;  /* CMP,L,A */
                {8'h61,8'h47,2'bxx} : dec_pc_inc2 = 1'b1;  /* CMP,H,A */
                {8'h4b,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* CMP,A,saddr */
                {8'h4e,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* CMP,A,[HL+byte] */
                {8'h61,8'hc0,2'bxx} : dec_pc_inc2 = 1'b1;  /* CMP,A,[HL+B] */
                {8'h61,8'hc2,2'bxx} : dec_pc_inc2 = 1'b1;  /* CMP,A,[HL+C] */
                {8'hd4,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* CMP0,,saddr */
                {8'h06,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDW,AX,saddrp */
                {8'h26,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBW,AX,saddrp */
                {8'h46,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* CMPW,AX,saddrp */
                {8'ha4,8'hxx,2'bx1} : dec_pc_inc2 = 1'b1;  /* INC,,saddr */
                {8'hb4,8'hxx,2'bx1} : dec_pc_inc2 = 1'b1;  /* DEC,,saddr */
                {8'ha6,8'hxx,2'bx1} : dec_pc_inc2 = 1'b1;  /* INCW,,saddrp */
                {8'hb6,8'hxx,2'bx1} : dec_pc_inc2 = 1'b1;  /* DECW,,saddrp */
                {8'h31,8'h0a,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHR,A,0 */
                {8'h31,8'h1a,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHR,A,1 */
                {8'h31,8'h2a,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHR,A,2 */
                {8'h31,8'h3a,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHR,A,3 */
                {8'h31,8'h4a,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHR,A,4 */
                {8'h31,8'h5a,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHR,A,5 */
                {8'h31,8'h6a,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHR,A,6 */
                {8'h31,8'h7a,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHR,A,7 */
                {8'h31,8'h0e,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,0 */
                {8'h31,8'h1e,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,1 */
                {8'h31,8'h2e,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,2 */
                {8'h31,8'h3e,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,3 */
                {8'h31,8'h4e,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,4 */
                {8'h31,8'h5e,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,5 */
                {8'h31,8'h6e,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,6 */
                {8'h31,8'h7e,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,7 */
                {8'h31,8'h8e,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,8 */
                {8'h31,8'h9e,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,9 */
                {8'h31,8'hae,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,10 */
                {8'h31,8'hbe,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,11 */
                {8'h31,8'hce,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,12 */
                {8'h31,8'hde,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,13 */
                {8'h31,8'hee,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,14 */
                {8'h31,8'hfe,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHRW,AX,15 */
                {8'h31,8'h09,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,A,0 */
                {8'h31,8'h19,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,A,1 */
                {8'h31,8'h29,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,A,2 */
                {8'h31,8'h39,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,A,3 */
                {8'h31,8'h49,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,A,4 */
                {8'h31,8'h59,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,A,5 */
                {8'h31,8'h69,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,A,6 */
                {8'h31,8'h79,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,A,7 */
                {8'h31,8'h08,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,B,0 */
                {8'h31,8'h18,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,B,1 */
                {8'h31,8'h28,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,B,2 */
                {8'h31,8'h38,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,B,3 */
                {8'h31,8'h48,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,B,4 */
                {8'h31,8'h58,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,B,5 */
                {8'h31,8'h68,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,B,6 */
                {8'h31,8'h78,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,B,7 */
                {8'h31,8'h07,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,C,0 */
                {8'h31,8'h17,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,C,1 */
                {8'h31,8'h27,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,C,2 */
                {8'h31,8'h37,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,C,3 */
                {8'h31,8'h47,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,C,4 */
                {8'h31,8'h57,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,C,5 */
                {8'h31,8'h67,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,C,6 */
                {8'h31,8'h77,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,C,7 */
                {8'h31,8'h0d,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,0 */
                {8'h31,8'h1d,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,1 */
                {8'h31,8'h2d,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,2 */
                {8'h31,8'h3d,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,3 */
                {8'h31,8'h4d,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,4 */
                {8'h31,8'h5d,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,5 */
                {8'h31,8'h6d,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,6 */
                {8'h31,8'h7d,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,7 */
                {8'h31,8'h8d,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,8 */
                {8'h31,8'h9d,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,9 */
                {8'h31,8'had,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,10 */
                {8'h31,8'hbd,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,11 */
                {8'h31,8'hcd,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,12 */
                {8'h31,8'hdd,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,13 */
                {8'h31,8'hed,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,14 */
                {8'h31,8'hfd,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,AX,15 */
                {8'h31,8'h0c,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,0 */
                {8'h31,8'h1c,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,1 */
                {8'h31,8'h2c,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,2 */
                {8'h31,8'h3c,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,3 */
                {8'h31,8'h4c,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,4 */
                {8'h31,8'h5c,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,5 */
                {8'h31,8'h6c,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,6 */
                {8'h31,8'h7c,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,7 */
                {8'h31,8'h8c,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,8 */
                {8'h31,8'h9c,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,9 */
                {8'h31,8'hac,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,10 */
                {8'h31,8'hbc,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,11 */
                {8'h31,8'hcc,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,12 */
                {8'h31,8'hdc,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,13 */
                {8'h31,8'hec,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,14 */
                {8'h31,8'hfc,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHLW,BC,15 */
                {8'h31,8'h0b,2'bxx} : dec_pc_inc2 = 1'b1;  /* SAR,A,0 */
                {8'h31,8'h1b,2'bxx} : dec_pc_inc2 = 1'b1;  /* SAR,A,1 */
                {8'h31,8'h2b,2'bxx} : dec_pc_inc2 = 1'b1;  /* SAR,A,2 */
                {8'h31,8'h3b,2'bxx} : dec_pc_inc2 = 1'b1;  /* SAR,A,3 */
                {8'h31,8'h4b,2'bxx} : dec_pc_inc2 = 1'b1;  /* SAR,A,4 */
                {8'h31,8'h5b,2'bxx} : dec_pc_inc2 = 1'b1;  /* SAR,A,5 */
                {8'h31,8'h6b,2'bxx} : dec_pc_inc2 = 1'b1;  /* SAR,A,6 */
                {8'h31,8'h7b,2'bxx} : dec_pc_inc2 = 1'b1;  /* SAR,A,7 */
                {8'h31,8'h0f,2'bxx} : dec_pc_inc2 = 1'b1;  /* SARW,AX,0 */
                {8'h31,8'h1f,2'bxx} : dec_pc_inc2 = 1'b1;  /* SARW,AX,1 */
                {8'h31,8'h2f,2'bxx} : dec_pc_inc2 = 1'b1;  /* SARW,AX,2 */
                {8'h31,8'h3f,2'bxx} : dec_pc_inc2 = 1'b1;  /* SARW,AX,3 */
                {8'h31,8'h4f,2'bxx} : dec_pc_inc2 = 1'b1;  /* SARW,AX,4 */
                {8'h31,8'h5f,2'bxx} : dec_pc_inc2 = 1'b1;  /* SARW,AX,5 */
                {8'h31,8'h6f,2'bxx} : dec_pc_inc2 = 1'b1;  /* SARW,AX,6 */
                {8'h31,8'h7f,2'bxx} : dec_pc_inc2 = 1'b1;  /* SARW,AX,7 */
                {8'h31,8'h8f,2'bxx} : dec_pc_inc2 = 1'b1;  /* SARW,AX,8 */
                {8'h31,8'h9f,2'bxx} : dec_pc_inc2 = 1'b1;  /* SARW,AX,9 */
                {8'h31,8'haf,2'bxx} : dec_pc_inc2 = 1'b1;  /* SARW,AX,10 */
                {8'h31,8'hbf,2'bxx} : dec_pc_inc2 = 1'b1;  /* SARW,AX,11 */
                {8'h31,8'hcf,2'bxx} : dec_pc_inc2 = 1'b1;  /* SARW,AX,12 */
                {8'h31,8'hdf,2'bxx} : dec_pc_inc2 = 1'b1;  /* SARW,AX,13 */
                {8'h31,8'hef,2'bxx} : dec_pc_inc2 = 1'b1;  /* SARW,AX,14 */
                {8'h31,8'hff,2'bxx} : dec_pc_inc2 = 1'b1;  /* SARW,AX,15 */
                {8'h61,8'hdb,2'bxx} : dec_pc_inc2 = 1'b1;  /* ROR,A,1 */
                {8'h61,8'heb,2'bxx} : dec_pc_inc2 = 1'b1;  /* ROL,A,1 */
                {8'h61,8'hfb,2'bxx} : dec_pc_inc2 = 1'b1;  /* RORC,A,1 */
                {8'h61,8'hdc,2'bxx} : dec_pc_inc2 = 1'b1;  /* ROLC,A,1 */
                {8'h61,8'hee,2'bxx} : dec_pc_inc2 = 1'b1;  /* ROLWC,AX,1 */
                {8'h61,8'hfe,2'bxx} : dec_pc_inc2 = 1'b1;  /* ROLWC,BC,1 */
                {8'h71,8'h8c,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,A.0 */
                {8'h71,8'h9c,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,A.1 */
                {8'h71,8'hac,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,A.2 */
                {8'h71,8'hbc,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,A.3 */
                {8'h71,8'hcc,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,A.4 */
                {8'h71,8'hdc,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,A.5 */
                {8'h71,8'hec,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,A.6 */
                {8'h71,8'hfc,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,A.7 */
                {8'h71,8'h84,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,[HL].0 */
                {8'h71,8'h94,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,[HL].1 */
                {8'h71,8'ha4,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,[HL].2 */
                {8'h71,8'hb4,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,[HL].3 */
                {8'h71,8'hc4,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,[HL].4 */
                {8'h71,8'hd4,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,[HL].5 */
                {8'h71,8'he4,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,[HL].6 */
                {8'h71,8'hf4,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,CY,[HL].7 */
                {8'h71,8'h89,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,A.0,CY */
                {8'h71,8'h99,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,A.1,CY */
                {8'h71,8'ha9,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,A.2,CY */
                {8'h71,8'hb9,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,A.3,CY */
                {8'h71,8'hc9,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,A.4,CY */
                {8'h71,8'hd9,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,A.5,CY */
                {8'h71,8'he9,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,A.6,CY */
                {8'h71,8'hf9,2'bxx} : dec_pc_inc2 = 1'b1;  /* MOV1,A.7,CY */
                {8'h71,8'h81,2'bx1} : dec_pc_inc2 = 1'b1;  /* MOV1,[HL].0,CY */
                {8'h71,8'h91,2'bx1} : dec_pc_inc2 = 1'b1;  /* MOV1,[HL].1,CY */
                {8'h71,8'ha1,2'bx1} : dec_pc_inc2 = 1'b1;  /* MOV1,[HL].2,CY */
                {8'h71,8'hb1,2'bx1} : dec_pc_inc2 = 1'b1;  /* MOV1,[HL].3,CY */
                {8'h71,8'hc1,2'bx1} : dec_pc_inc2 = 1'b1;  /* MOV1,[HL].4,CY */
                {8'h71,8'hd1,2'bx1} : dec_pc_inc2 = 1'b1;  /* MOV1,[HL].5,CY */
                {8'h71,8'he1,2'bx1} : dec_pc_inc2 = 1'b1;  /* MOV1,[HL].6,CY */
                {8'h71,8'hf1,2'bx1} : dec_pc_inc2 = 1'b1;  /* MOV1,[HL].7,CY */
                {8'h71,8'h8d,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND1,CY,A.0 */
                {8'h71,8'h9d,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND1,CY,A.1 */
                {8'h71,8'had,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND1,CY,A.2 */
                {8'h71,8'hbd,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND1,CY,A.3 */
                {8'h71,8'hcd,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND1,CY,A.4 */
                {8'h71,8'hdd,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND1,CY,A.5 */
                {8'h71,8'hed,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND1,CY,A.6 */
                {8'h71,8'hfd,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND1,CY,A.7 */
                {8'h71,8'h85,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND1,CY,[HL].0 */
                {8'h71,8'h95,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND1,CY,[HL].1 */
                {8'h71,8'ha5,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND1,CY,[HL].2 */
                {8'h71,8'hb5,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND1,CY,[HL].3 */
                {8'h71,8'hc5,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND1,CY,[HL].4 */
                {8'h71,8'hd5,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND1,CY,[HL].5 */
                {8'h71,8'he5,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND1,CY,[HL].6 */
                {8'h71,8'hf5,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND1,CY,[HL].7 */
                {8'h71,8'h8e,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR1,CY,A.0 */
                {8'h71,8'h9e,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR1,CY,A.1 */
                {8'h71,8'hae,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR1,CY,A.2 */
                {8'h71,8'hbe,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR1,CY,A.3 */
                {8'h71,8'hce,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR1,CY,A.4 */
                {8'h71,8'hde,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR1,CY,A.5 */
                {8'h71,8'hee,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR1,CY,A.6 */
                {8'h71,8'hfe,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR1,CY,A.7 */
                {8'h71,8'h86,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR1,CY,[HL].0 */
                {8'h71,8'h96,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR1,CY,[HL].1 */
                {8'h71,8'ha6,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR1,CY,[HL].2 */
                {8'h71,8'hb6,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR1,CY,[HL].3 */
                {8'h71,8'hc6,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR1,CY,[HL].4 */
                {8'h71,8'hd6,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR1,CY,[HL].5 */
                {8'h71,8'he6,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR1,CY,[HL].6 */
                {8'h71,8'hf6,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR1,CY,[HL].7 */
                {8'h71,8'h8f,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,A.0 */
                {8'h71,8'h9f,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,A.1 */
                {8'h71,8'haf,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,A.2 */
                {8'h71,8'hbf,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,A.3 */
                {8'h71,8'hcf,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,A.4 */
                {8'h71,8'hdf,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,A.5 */
                {8'h71,8'hef,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,A.6 */
                {8'h71,8'hff,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,A.7 */
                {8'h71,8'h87,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,[HL].0 */
                {8'h71,8'h97,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,[HL].1 */
                {8'h71,8'ha7,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,[HL].2 */
                {8'h71,8'hb7,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,[HL].3 */
                {8'h71,8'hc7,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,[HL].4 */
                {8'h71,8'hd7,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,[HL].5 */
                {8'h71,8'he7,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,[HL].6 */
                {8'h71,8'hf7,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR1,CY,[HL].7 */
                {8'h71,8'h8a,2'bxx} : dec_pc_inc2 = 1'b1;  /* SET1,,A.0 */
                {8'h71,8'h9a,2'bxx} : dec_pc_inc2 = 1'b1;  /* SET1,,A.1 */
                {8'h71,8'haa,2'bxx} : dec_pc_inc2 = 1'b1;  /* SET1,,A.2 */
                {8'h71,8'hba,2'bxx} : dec_pc_inc2 = 1'b1;  /* SET1,,A.3 */
                {8'h71,8'hca,2'bxx} : dec_pc_inc2 = 1'b1;  /* SET1,,A.4 */
                {8'h71,8'hda,2'bxx} : dec_pc_inc2 = 1'b1;  /* SET1,,A.5 */
                {8'h71,8'hea,2'bxx} : dec_pc_inc2 = 1'b1;  /* SET1,,A.6 */
                {8'h71,8'hfa,2'bxx} : dec_pc_inc2 = 1'b1;  /* SET1,,A.7 */
                {8'h71,8'h82,2'bx1} : dec_pc_inc2 = 1'b1;  /* SET1,,[HL].0 */
                {8'h71,8'h92,2'bx1} : dec_pc_inc2 = 1'b1;  /* SET1,,[HL].1 */
                {8'h71,8'ha2,2'bx1} : dec_pc_inc2 = 1'b1;  /* SET1,,[HL].2 */
                {8'h71,8'hb2,2'bx1} : dec_pc_inc2 = 1'b1;  /* SET1,,[HL].3 */
                {8'h71,8'hc2,2'bx1} : dec_pc_inc2 = 1'b1;  /* SET1,,[HL].4 */
                {8'h71,8'hd2,2'bx1} : dec_pc_inc2 = 1'b1;  /* SET1,,[HL].5 */
                {8'h71,8'he2,2'bx1} : dec_pc_inc2 = 1'b1;  /* SET1,,[HL].6 */
                {8'h71,8'hf2,2'bx1} : dec_pc_inc2 = 1'b1;  /* SET1,,[HL].7 */
                {8'h71,8'h8b,2'bxx} : dec_pc_inc2 = 1'b1;  /* CLR1,,A.0 */
                {8'h71,8'h9b,2'bxx} : dec_pc_inc2 = 1'b1;  /* CLR1,,A.1 */
                {8'h71,8'hab,2'bxx} : dec_pc_inc2 = 1'b1;  /* CLR1,,A.2 */
                {8'h71,8'hbb,2'bxx} : dec_pc_inc2 = 1'b1;  /* CLR1,,A.3 */
                {8'h71,8'hcb,2'bxx} : dec_pc_inc2 = 1'b1;  /* CLR1,,A.4 */
                {8'h71,8'hdb,2'bxx} : dec_pc_inc2 = 1'b1;  /* CLR1,,A.5 */
                {8'h71,8'heb,2'bxx} : dec_pc_inc2 = 1'b1;  /* CLR1,,A.6 */
                {8'h71,8'hfb,2'bxx} : dec_pc_inc2 = 1'b1;  /* CLR1,,A.7 */
                {8'h71,8'h83,2'bx1} : dec_pc_inc2 = 1'b1;  /* CLR1,,[HL].0 */
                {8'h71,8'h93,2'bx1} : dec_pc_inc2 = 1'b1;  /* CLR1,,[HL].1 */
                {8'h71,8'ha3,2'bx1} : dec_pc_inc2 = 1'b1;  /* CLR1,,[HL].2 */
                {8'h71,8'hb3,2'bx1} : dec_pc_inc2 = 1'b1;  /* CLR1,,[HL].3 */
                {8'h71,8'hc3,2'bx1} : dec_pc_inc2 = 1'b1;  /* CLR1,,[HL].4 */
                {8'h71,8'hd3,2'bx1} : dec_pc_inc2 = 1'b1;  /* CLR1,,[HL].5 */
                {8'h71,8'he3,2'bx1} : dec_pc_inc2 = 1'b1;  /* CLR1,,[HL].6 */
                {8'h71,8'hf3,2'bx1} : dec_pc_inc2 = 1'b1;  /* CLR1,,[HL].7 */
                {8'h71,8'h80,2'bxx} : dec_pc_inc2 = 1'b1;  /* SET1,,CY */
                {8'h71,8'h88,2'bxx} : dec_pc_inc2 = 1'b1;  /* CLR1,,CY */
                {8'h71,8'hc0,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOT1,,CY */
                {8'h61,8'hca,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALL,,AX */
                {8'h61,8'hda,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALL,,BC */
                {8'h61,8'hea,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALL,,DE */
                {8'h61,8'hfa,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALL,,HL */
                {8'h61,8'h84,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[0080h] */
                {8'h61,8'h94,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[0082h] */
                {8'h61,8'ha4,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[0084h] */
                {8'h61,8'hb4,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[0086h] */
                {8'h61,8'hc4,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[0088h] */
                {8'h61,8'hd4,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[008Ah] */
                {8'h61,8'he4,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[008Ch] */
                {8'h61,8'hf4,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[008Eh] */
                {8'h61,8'h85,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[0090h] */
                {8'h61,8'h95,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[0092h] */
                {8'h61,8'ha5,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[0094h] */
                {8'h61,8'hb5,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[0096h] */
                {8'h61,8'hc5,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[0098h] */
                {8'h61,8'hd5,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[009Ah] */
                {8'h61,8'he5,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[009Ch] */
                {8'h61,8'hf5,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[009Eh] */
                {8'h61,8'h86,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00A0h] */
                {8'h61,8'h96,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00A2h] */
                {8'h61,8'ha6,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00A4h] */
                {8'h61,8'hb6,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00A6h] */
                {8'h61,8'hc6,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00A8h] */
                {8'h61,8'hd6,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00AAh] */
                {8'h61,8'he6,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00ACh] */
                {8'h61,8'hf6,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00AEh] */
                {8'h61,8'h87,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00B0h] */
                {8'h61,8'h97,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00B2h] */
                {8'h61,8'ha7,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00B4h] */
                {8'h61,8'hb7,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00B6h] */
                {8'h61,8'hc7,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00B8h] */
                {8'h61,8'hd7,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00BAh] */
                {8'h61,8'he7,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00BCh] */
                {8'h61,8'hf7,2'bx0} : dec_pc_inc2 = 1'b1;  /* CALLT,,[00BEh] */
                {8'h61,8'hcc,2'bx0} : dec_pc_inc2 = 1'b1;  /* BRK,, */
                {8'h61,8'hdd,2'bxx} : dec_pc_inc2 = 1'b1;  /* PUSH,,PSW */
                {8'h61,8'hcd,2'bxx} : dec_pc_inc2 = 1'b1;  /* POP,,PSW */
                {8'h10,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDW,SP,#byte */
                {8'h20,8'hxx,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBW,SP,#byte */
                {8'hef,8'hxx,2'bx0} : dec_pc_inc2 = 1'b1;  /* BR,,$addr8 */
                {8'h61,8'hcb,2'bx0} : dec_pc_inc2 = 1'b1;  /* BR,,AX */
                {8'hdc,8'hxx,2'bx1} : dec_pc_inc2 = 1'b1;  /* BC,,$addr8 */
                {8'hde,8'hxx,2'bx1} : dec_pc_inc2 = 1'b1;  /* BNC,,$addr8 */
                {8'hdd,8'hxx,2'bx1} : dec_pc_inc2 = 1'b1;  /* BZ,,$addr8 */
                {8'hdf,8'hxx,2'bx1} : dec_pc_inc2 = 1'b1;  /* BNZ,,$addr8 */
                {8'h61,8'hc8,2'bxx} : dec_pc_inc2 = 1'b1;  /* SKC,, */
                {8'h61,8'hd8,2'bxx} : dec_pc_inc2 = 1'b1;  /* SKNC,, */
                {8'h61,8'he8,2'bxx} : dec_pc_inc2 = 1'b1;  /* SKZ,, */
                {8'h61,8'hf8,2'bxx} : dec_pc_inc2 = 1'b1;  /* SKNZ,, */
                {8'h61,8'he3,2'bxx} : dec_pc_inc2 = 1'b1;  /* SKH,, */
                {8'h61,8'hf3,2'bxx} : dec_pc_inc2 = 1'b1;  /* SKNH,, */
                {8'h61,8'hcf,2'bxx} : dec_pc_inc2 = 1'b1;  /* SEL,,RB0 */
                {8'h61,8'hdf,2'bxx} : dec_pc_inc2 = 1'b1;  /* SEL,,RB1 */
                {8'h61,8'hef,2'bxx} : dec_pc_inc2 = 1'b1;  /* SEL,,RB2 */
                {8'h61,8'hff,2'bxx} : dec_pc_inc2 = 1'b1;  /* SEL,,RB3 */
                {8'h61,8'hed,2'b10} : dec_pc_inc2 = 1'b1;  /* HALT,, */
                {8'h61,8'hfd,2'b10} : dec_pc_inc2 = 1'b1;  /* STOP,, */
                {8'h61,8'ha1,2'bx0} : dec_pc_inc2 = 1'b1;  /* SOFT2,,BREAK */
                {8'h61,8'h81,2'bxx} : dec_pc_inc2 = 1'b1;  /* ALT1,, */
                {8'h61,8'h91,2'bxx} : dec_pc_inc2 = 1'b1;  /* ALT2,, */
                {8'h61,8'h88,2'bxx} : dec_pc_inc2 = 1'b1;  /* XCH,A,X */
                {8'h61,8'h98,2'bxx} : dec_pc_inc2 = 1'b1;  /* XCH,A,X */
                {8'h61,8'h99,2'bxx} : dec_pc_inc2 = 1'b1;  /* XCH,A,X */
                {8'h61,8'h9a,2'bxx} : dec_pc_inc2 = 1'b1;  /* XCH,A,C */
                {8'h61,8'h9b,2'bxx} : dec_pc_inc2 = 1'b1;  /* XCH,A,B */
                {8'h61,8'h9c,2'bxx} : dec_pc_inc2 = 1'b1;  /* XCH,A,E */
                {8'h61,8'h9d,2'bxx} : dec_pc_inc2 = 1'b1;  /* XCH,A,D */
                {8'h61,8'h9e,2'bxx} : dec_pc_inc2 = 1'b1;  /* XCH,A,L */
                {8'h61,8'h9f,2'bxx} : dec_pc_inc2 = 1'b1;  /* XCH,A,H */
                {8'h61,8'hbe,2'bx1} : dec_pc_inc2 = 1'b1;  /* XCH,A,[DE] */
                {8'h61,8'hbc,2'bx1} : dec_pc_inc2 = 1'b1;  /* XCH,A,[HL] */
                {8'h61,8'h19,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDC,A,A */
                {8'h61,8'h39,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBC,A,A */
                {8'h61,8'hd1,2'bxx} : dec_pc_inc2 = 1'b1;  /* AND,A,[HL+B] */
                {8'h61,8'he1,2'bxx} : dec_pc_inc2 = 1'b1;  /* OR,A,[HL+B] */
                {8'h61,8'hf1,2'bxx} : dec_pc_inc2 = 1'b1;  /* XOR,A,[HL+B] */
                {8'h61,8'h83,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADD,A,[HL+C] */
                {8'h61,8'h93,2'bxx} : dec_pc_inc2 = 1'b1;  /* ADDC,A,[HL+C] */
                {8'h61,8'ha3,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUB,A,[HL+C] */
                {8'h61,8'hb3,2'bxx} : dec_pc_inc2 = 1'b1;  /* SUBC,A,[HL+C] */
                {8'h71,8'h90,2'bxx} : dec_pc_inc2 = 1'b1;  /* SET1,,CY */
                {8'h71,8'ha0,2'bxx} : dec_pc_inc2 = 1'b1;  /* SET1,,CY */
                {8'h71,8'hb0,2'bxx} : dec_pc_inc2 = 1'b1;  /* SET1,,CY */
                {8'h71,8'hd0,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOT1,,CY */
                {8'h71,8'he0,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOT1,,CY */
                {8'h71,8'hf0,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOT1,,CY */
                {8'h71,8'h98,2'bxx} : dec_pc_inc2 = 1'b1;  /* CLR1,,CY */
                {8'h71,8'ha8,2'bxx} : dec_pc_inc2 = 1'b1;  /* CLR1,,CY */
                {8'h71,8'hb8,2'bxx} : dec_pc_inc2 = 1'b1;  /* CLR1,,CY */
                {8'h71,8'hc8,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOT1,,CY */
                {8'h71,8'hd8,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOT1,,CY */
                {8'h71,8'he8,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOT1,,CY */
                {8'h71,8'hf8,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOT1,,CY */
                {8'h31,8'h8a,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHR,A,0 */
                {8'h31,8'h9a,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHR,A,1 */
                {8'h31,8'haa,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHR,A,2 */
                {8'h31,8'hba,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHR,A,3 */
                {8'h31,8'hca,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHR,A,4 */
                {8'h31,8'hda,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHR,A,5 */
                {8'h31,8'hea,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHR,A,6 */
                {8'h31,8'hfa,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHR,A,7 */
                {8'h31,8'h89,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,A,0 */
                {8'h31,8'h99,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,A,1 */
                {8'h31,8'ha9,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,A,2 */
                {8'h31,8'hb9,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,A,3 */
                {8'h31,8'hc9,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,A,4 */
                {8'h31,8'hd9,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,A,5 */
                {8'h31,8'he9,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,A,6 */
                {8'h31,8'hf9,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,A,7 */
                {8'h31,8'h88,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,B,0 */
                {8'h31,8'h98,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,B,1 */
                {8'h31,8'ha8,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,B,2 */
                {8'h31,8'hb8,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,B,3 */
                {8'h31,8'hc8,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,B,4 */
                {8'h31,8'hd8,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,B,5 */
                {8'h31,8'he8,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,B,6 */
                {8'h31,8'hf8,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,B,7 */
                {8'h31,8'h87,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,C,0 */
                {8'h31,8'h97,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,C,1 */
                {8'h31,8'ha7,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,C,2 */
                {8'h31,8'hb7,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,C,3 */
                {8'h31,8'hc7,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,C,4 */
                {8'h31,8'hd7,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,C,5 */
                {8'h31,8'he7,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,C,6 */
                {8'h31,8'hf7,2'bxx} : dec_pc_inc2 = 1'b1;  /* SHL,C,7 */
                {8'h31,8'h8b,2'bxx} : dec_pc_inc2 = 1'b1;  /* SAR,A,0 */
                {8'h31,8'h9b,2'bxx} : dec_pc_inc2 = 1'b1;  /* SAR,A,1 */
                {8'h31,8'hab,2'bxx} : dec_pc_inc2 = 1'b1;  /* SAR,A,2 */
                {8'h31,8'hbb,2'bxx} : dec_pc_inc2 = 1'b1;  /* SAR,A,3 */
                {8'h31,8'hcb,2'bxx} : dec_pc_inc2 = 1'b1;  /* SAR,A,4 */
                {8'h31,8'hdb,2'bxx} : dec_pc_inc2 = 1'b1;  /* SAR,A,5 */
                {8'h31,8'heb,2'bxx} : dec_pc_inc2 = 1'b1;  /* SAR,A,6 */
                {8'h31,8'hfb,2'bxx} : dec_pc_inc2 = 1'b1;  /* SAR,A,7 */
                {8'h31,8'h06,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'h16,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'h26,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'h36,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'h46,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'h56,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'h66,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'h76,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'h86,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'h96,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'ha6,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'hb6,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'hc6,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'hd6,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'he6,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                {8'h31,8'hf6,2'bxx} : dec_pc_inc2 = 1'b1;  /* NOP,, */
                default : dec_pc_inc2 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_pc_inc3;
    reg    dec_pc_inc3;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1) begin
            dec_pc_inc3 = 1'b0;
        end else if(skpack == 1'b1) begin
            casex ({ID_stage0,ID_stage1})  
                {8'hcd,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOV,saddr,#byte */
                {8'hce,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOV,sfr,#byte */
                {8'hca,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOV,[DE+byte],#byte */
                {8'hcc,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOV,[HL+byte],#byte */
                {8'h8f,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOV,A,!addr16 */
                {8'h9f,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOV,!addr16,A */
                {8'h09,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOV,A,word[B] */
                {8'h18,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOV,word[B],A */
                {8'h29,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOV,A,word[C] */
                {8'h28,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOV,word[C],A */
                {8'h49,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOV,A,word[BC] */
                {8'h48,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOV,word[BC],A */
                {8'hc8,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOV,[SP+byte],#byte */
                {8'he9,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOV,B,!addr16 */
                {8'hf9,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOV,C,!addr16 */
                {8'hd9,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOV,X,!addr16 */
                {8'h61,8'hb8} : dec_pc_inc3 = 1'b1;  /* MOV,ES,saddr */
                {8'h61,8'hce} : dec_pc_inc3 = 1'b1;  /* MOVS,[HL+byte],X */
                {8'h61,8'ha8} : dec_pc_inc3 = 1'b1;  /* XCH,A,saddr */
                {8'h61,8'hab} : dec_pc_inc3 = 1'b1;  /* XCH,A,sfr */
                {8'h61,8'haf} : dec_pc_inc3 = 1'b1;  /* XCH,A,[DE+byte] */
                {8'h61,8'had} : dec_pc_inc3 = 1'b1;  /* XCH,A,[HL+byte] */
                {8'he5,8'hxx} : dec_pc_inc3 = 1'b1;  /* ONEB,,!addr16 */
                {8'hf5,8'hxx} : dec_pc_inc3 = 1'b1;  /* CLRB,,!addr16 */
                {8'h30,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOVW,AX,#word */
                {8'h32,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOVW,BC,#word */
                {8'h34,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOVW,DE,#word */
                {8'h36,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOVW,HL,#word */
                {8'haf,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOVW,AX,!addr16 */
                {8'hbf,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOVW,!addr16,AX */
                {8'h59,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOVW,AX,word[B] */
                {8'h58,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOVW,word[B],AX */
                {8'h69,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOVW,AX,word[C] */
                {8'h68,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOVW,word[C],AX */
                {8'h79,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOVW,AX,word[BC] */
                {8'h78,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOVW,word[BC],AX */
                {8'hdb,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOVW,BC,!addr16 */
                {8'heb,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOVW,DE,!addr16 */
                {8'hfb,8'hxx} : dec_pc_inc3 = 1'b1;  /* MOVW,HL,!addr16 */
                {8'h0a,8'hxx} : dec_pc_inc3 = 1'b1;  /* ADD,saddr,#byte */
                {8'h0f,8'hxx} : dec_pc_inc3 = 1'b1;  /* ADD,A,!addr16 */
                {8'h1a,8'hxx} : dec_pc_inc3 = 1'b1;  /* ADDC,saddr,#byte */
                {8'h1f,8'hxx} : dec_pc_inc3 = 1'b1;  /* ADDC,A,!addr16 */
                {8'h2a,8'hxx} : dec_pc_inc3 = 1'b1;  /* SUB,saddr,#byte */
                {8'h2f,8'hxx} : dec_pc_inc3 = 1'b1;  /* SUB,A,!addr16 */
                {8'h3a,8'hxx} : dec_pc_inc3 = 1'b1;  /* SUBC,saddr,#byte */
                {8'h3f,8'hxx} : dec_pc_inc3 = 1'b1;  /* SUBC,A,!addr16 */
                {8'h5a,8'hxx} : dec_pc_inc3 = 1'b1;  /* AND,saddr,#byte */
                {8'h5f,8'hxx} : dec_pc_inc3 = 1'b1;  /* AND,A,!addr16 */
                {8'h6a,8'hxx} : dec_pc_inc3 = 1'b1;  /* OR,saddr,#byte */
                {8'h6f,8'hxx} : dec_pc_inc3 = 1'b1;  /* OR,A,!addr16 */
                {8'h7a,8'hxx} : dec_pc_inc3 = 1'b1;  /* XOR,saddr,#byte */
                {8'h7f,8'hxx} : dec_pc_inc3 = 1'b1;  /* XOR,A,!addr16 */
                {8'h4a,8'hxx} : dec_pc_inc3 = 1'b1;  /* CMP,saddr,#byte */
                {8'h4f,8'hxx} : dec_pc_inc3 = 1'b1;  /* CMP,A,!addr16 */
                {8'h61,8'hde} : dec_pc_inc3 = 1'b1;  /* CMPS,X,[HL+byte] */
                {8'hd5,8'hxx} : dec_pc_inc3 = 1'b1;  /* CMP0,,!addr16 */
                {8'h04,8'hxx} : dec_pc_inc3 = 1'b1;  /* ADDW,AX,#word */
                {8'h02,8'hxx} : dec_pc_inc3 = 1'b1;  /* ADDW,AX,!addr16 */
                {8'h61,8'h09} : dec_pc_inc3 = 1'b1;  /* ADDW,AX,[HL+byte] */
                {8'h24,8'hxx} : dec_pc_inc3 = 1'b1;  /* SUBW,AX,#word */
                {8'h22,8'hxx} : dec_pc_inc3 = 1'b1;  /* SUBW,AX,!addr16 */
                {8'h61,8'h29} : dec_pc_inc3 = 1'b1;  /* SUBW,AX,[HL+byte] */
                {8'h44,8'hxx} : dec_pc_inc3 = 1'b1;  /* CMPW,AX,#word */
                {8'h42,8'hxx} : dec_pc_inc3 = 1'b1;  /* CMPW,AX,!addr16 */
                {8'h61,8'h49} : dec_pc_inc3 = 1'b1;  /* CMPW,AX,[HL+byte] */
                {8'ha0,8'hxx} : dec_pc_inc3 = 1'b1;  /* INC,,!addr16 */
                {8'h61,8'h59} : dec_pc_inc3 = 1'b1;  /* INC,,[HL+byte] */
                {8'hb0,8'hxx} : dec_pc_inc3 = 1'b1;  /* DEC,,!addr16 */
                {8'h61,8'h69} : dec_pc_inc3 = 1'b1;  /* DEC,,[HL+byte] */
                {8'ha2,8'hxx} : dec_pc_inc3 = 1'b1;  /* INCW,,!addr16 */
                {8'h61,8'h79} : dec_pc_inc3 = 1'b1;  /* INCW,,[HL+byte] */
                {8'hb2,8'hxx} : dec_pc_inc3 = 1'b1;  /* DECW,,!addr16 */
                {8'h61,8'h89} : dec_pc_inc3 = 1'b1;  /* DECW,,[HL+byte] */
                {8'h71,8'h04} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,saddr.0 */
                {8'h71,8'h14} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,saddr.1 */
                {8'h71,8'h24} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,saddr.2 */
                {8'h71,8'h34} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,saddr.3 */
                {8'h71,8'h44} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,saddr.4 */
                {8'h71,8'h54} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,saddr.5 */
                {8'h71,8'h64} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,saddr.6 */
                {8'h71,8'h74} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,saddr.7 */
                {8'h71,8'h0c} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,sfr.0 */
                {8'h71,8'h1c} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,sfr.1 */
                {8'h71,8'h2c} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,sfr.2 */
                {8'h71,8'h3c} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,sfr.3 */
                {8'h71,8'h4c} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,sfr.4 */
                {8'h71,8'h5c} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,sfr.5 */
                {8'h71,8'h6c} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,sfr.6 */
                {8'h71,8'h7c} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,sfr.7 */
                {8'h71,8'h01} : dec_pc_inc3 = 1'b1;  /* MOV1,saddr.0,CY */
                {8'h71,8'h11} : dec_pc_inc3 = 1'b1;  /* MOV1,saddr.1,CY */
                {8'h71,8'h21} : dec_pc_inc3 = 1'b1;  /* MOV1,saddr.2,CY */
                {8'h71,8'h31} : dec_pc_inc3 = 1'b1;  /* MOV1,saddr.3,CY */
                {8'h71,8'h41} : dec_pc_inc3 = 1'b1;  /* MOV1,saddr.4,CY */
                {8'h71,8'h51} : dec_pc_inc3 = 1'b1;  /* MOV1,saddr.5,CY */
                {8'h71,8'h61} : dec_pc_inc3 = 1'b1;  /* MOV1,saddr.6,CY */
                {8'h71,8'h71} : dec_pc_inc3 = 1'b1;  /* MOV1,saddr.7,CY */
                {8'h71,8'h09} : dec_pc_inc3 = 1'b1;  /* MOV1,sfr.0,CY */
                {8'h71,8'h19} : dec_pc_inc3 = 1'b1;  /* MOV1,sfr.1,CY */
                {8'h71,8'h29} : dec_pc_inc3 = 1'b1;  /* MOV1,sfr.2,CY */
                {8'h71,8'h39} : dec_pc_inc3 = 1'b1;  /* MOV1,sfr.3,CY */
                {8'h71,8'h49} : dec_pc_inc3 = 1'b1;  /* MOV1,sfr.4,CY */
                {8'h71,8'h59} : dec_pc_inc3 = 1'b1;  /* MOV1,sfr.5,CY */
                {8'h71,8'h69} : dec_pc_inc3 = 1'b1;  /* MOV1,sfr.6,CY */
                {8'h71,8'h79} : dec_pc_inc3 = 1'b1;  /* MOV1,sfr.7,CY */
                {8'h71,8'h05} : dec_pc_inc3 = 1'b1;  /* AND1,CY,saddr.0 */
                {8'h71,8'h15} : dec_pc_inc3 = 1'b1;  /* AND1,CY,saddr.1 */
                {8'h71,8'h25} : dec_pc_inc3 = 1'b1;  /* AND1,CY,saddr.2 */
                {8'h71,8'h35} : dec_pc_inc3 = 1'b1;  /* AND1,CY,saddr.3 */
                {8'h71,8'h45} : dec_pc_inc3 = 1'b1;  /* AND1,CY,saddr.4 */
                {8'h71,8'h55} : dec_pc_inc3 = 1'b1;  /* AND1,CY,saddr.5 */
                {8'h71,8'h65} : dec_pc_inc3 = 1'b1;  /* AND1,CY,saddr.6 */
                {8'h71,8'h75} : dec_pc_inc3 = 1'b1;  /* AND1,CY,saddr.7 */
                {8'h71,8'h0d} : dec_pc_inc3 = 1'b1;  /* AND1,CY,sfr.0 */
                {8'h71,8'h1d} : dec_pc_inc3 = 1'b1;  /* AND1,CY,sfr.1 */
                {8'h71,8'h2d} : dec_pc_inc3 = 1'b1;  /* AND1,CY,sfr.2 */
                {8'h71,8'h3d} : dec_pc_inc3 = 1'b1;  /* AND1,CY,sfr.3 */
                {8'h71,8'h4d} : dec_pc_inc3 = 1'b1;  /* AND1,CY,sfr.4 */
                {8'h71,8'h5d} : dec_pc_inc3 = 1'b1;  /* AND1,CY,sfr.5 */
                {8'h71,8'h6d} : dec_pc_inc3 = 1'b1;  /* AND1,CY,sfr.6 */
                {8'h71,8'h7d} : dec_pc_inc3 = 1'b1;  /* AND1,CY,sfr.7 */
                {8'h71,8'h06} : dec_pc_inc3 = 1'b1;  /* OR1,CY,saddr.0 */
                {8'h71,8'h16} : dec_pc_inc3 = 1'b1;  /* OR1,CY,saddr.1 */
                {8'h71,8'h26} : dec_pc_inc3 = 1'b1;  /* OR1,CY,saddr.2 */
                {8'h71,8'h36} : dec_pc_inc3 = 1'b1;  /* OR1,CY,saddr.3 */
                {8'h71,8'h46} : dec_pc_inc3 = 1'b1;  /* OR1,CY,saddr.4 */
                {8'h71,8'h56} : dec_pc_inc3 = 1'b1;  /* OR1,CY,saddr.5 */
                {8'h71,8'h66} : dec_pc_inc3 = 1'b1;  /* OR1,CY,saddr.6 */
                {8'h71,8'h76} : dec_pc_inc3 = 1'b1;  /* OR1,CY,saddr.7 */
                {8'h71,8'h0e} : dec_pc_inc3 = 1'b1;  /* OR1,CY,sfr.0 */
                {8'h71,8'h1e} : dec_pc_inc3 = 1'b1;  /* OR1,CY,sfr.1 */
                {8'h71,8'h2e} : dec_pc_inc3 = 1'b1;  /* OR1,CY,sfr.2 */
                {8'h71,8'h3e} : dec_pc_inc3 = 1'b1;  /* OR1,CY,sfr.3 */
                {8'h71,8'h4e} : dec_pc_inc3 = 1'b1;  /* OR1,CY,sfr.4 */
                {8'h71,8'h5e} : dec_pc_inc3 = 1'b1;  /* OR1,CY,sfr.5 */
                {8'h71,8'h6e} : dec_pc_inc3 = 1'b1;  /* OR1,CY,sfr.6 */
                {8'h71,8'h7e} : dec_pc_inc3 = 1'b1;  /* OR1,CY,sfr.7 */
                {8'h71,8'h07} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,saddr.0 */
                {8'h71,8'h17} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,saddr.1 */
                {8'h71,8'h27} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,saddr.2 */
                {8'h71,8'h37} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,saddr.3 */
                {8'h71,8'h47} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,saddr.4 */
                {8'h71,8'h57} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,saddr.5 */
                {8'h71,8'h67} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,saddr.6 */
                {8'h71,8'h77} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,saddr.7 */
                {8'h71,8'h0f} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,sfr.0 */
                {8'h71,8'h1f} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,sfr.1 */
                {8'h71,8'h2f} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,sfr.2 */
                {8'h71,8'h3f} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,sfr.3 */
                {8'h71,8'h4f} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,sfr.4 */
                {8'h71,8'h5f} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,sfr.5 */
                {8'h71,8'h6f} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,sfr.6 */
                {8'h71,8'h7f} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,sfr.7 */
                {8'h71,8'h02} : dec_pc_inc3 = 1'b1;  /* SET1,,saddr.0 */
                {8'h71,8'h12} : dec_pc_inc3 = 1'b1;  /* SET1,,saddr.1 */
                {8'h71,8'h22} : dec_pc_inc3 = 1'b1;  /* SET1,,saddr.2 */
                {8'h71,8'h32} : dec_pc_inc3 = 1'b1;  /* SET1,,saddr.3 */
                {8'h71,8'h42} : dec_pc_inc3 = 1'b1;  /* SET1,,saddr.4 */
                {8'h71,8'h52} : dec_pc_inc3 = 1'b1;  /* SET1,,saddr.5 */
                {8'h71,8'h62} : dec_pc_inc3 = 1'b1;  /* SET1,,saddr.6 */
                {8'h71,8'h72} : dec_pc_inc3 = 1'b1;  /* SET1,,saddr.7 */
                {8'h71,8'h0a} : dec_pc_inc3 = 1'b1;  /* SET1,,sfr.0 */
                {8'h71,8'h1a} : dec_pc_inc3 = 1'b1;  /* SET1,,sfr.1 */
                {8'h71,8'h2a} : dec_pc_inc3 = 1'b1;  /* SET1,,sfr.2 */
                {8'h71,8'h3a} : dec_pc_inc3 = 1'b1;  /* SET1,,sfr.3 */
                {8'h71,8'h4a} : dec_pc_inc3 = 1'b1;  /* SET1,,sfr.4 */
                {8'h71,8'h5a} : dec_pc_inc3 = 1'b1;  /* SET1,,sfr.5 */
                {8'h71,8'h6a} : dec_pc_inc3 = 1'b1;  /* SET1,,sfr.6 */
                {8'h71,8'h7a} : dec_pc_inc3 = 1'b1;  /* SET1,,sfr.7 */
                {8'h71,8'h03} : dec_pc_inc3 = 1'b1;  /* CLR1,,saddr.0 */
                {8'h71,8'h13} : dec_pc_inc3 = 1'b1;  /* CLR1,,saddr.1 */
                {8'h71,8'h23} : dec_pc_inc3 = 1'b1;  /* CLR1,,saddr.2 */
                {8'h71,8'h33} : dec_pc_inc3 = 1'b1;  /* CLR1,,saddr.3 */
                {8'h71,8'h43} : dec_pc_inc3 = 1'b1;  /* CLR1,,saddr.4 */
                {8'h71,8'h53} : dec_pc_inc3 = 1'b1;  /* CLR1,,saddr.5 */
                {8'h71,8'h63} : dec_pc_inc3 = 1'b1;  /* CLR1,,saddr.6 */
                {8'h71,8'h73} : dec_pc_inc3 = 1'b1;  /* CLR1,,saddr.7 */
                {8'h71,8'h0b} : dec_pc_inc3 = 1'b1;  /* CLR1,,sfr.0 */
                {8'h71,8'h1b} : dec_pc_inc3 = 1'b1;  /* CLR1,,sfr.1 */
                {8'h71,8'h2b} : dec_pc_inc3 = 1'b1;  /* CLR1,,sfr.2 */
                {8'h71,8'h3b} : dec_pc_inc3 = 1'b1;  /* CLR1,,sfr.3 */
                {8'h71,8'h4b} : dec_pc_inc3 = 1'b1;  /* CLR1,,sfr.4 */
                {8'h71,8'h5b} : dec_pc_inc3 = 1'b1;  /* CLR1,,sfr.5 */
                {8'h71,8'h6b} : dec_pc_inc3 = 1'b1;  /* CLR1,,sfr.6 */
                {8'h71,8'h7b} : dec_pc_inc3 = 1'b1;  /* CLR1,,sfr.7 */
                {8'hfe,8'hxx} : dec_pc_inc3 = 1'b1;  /* CALL,,$!addr16 */
                {8'hfd,8'hxx} : dec_pc_inc3 = 1'b1;  /* CALL,,!addr16 */
                {8'hed,8'hxx} : dec_pc_inc3 = 1'b1;  /* BR,,!addr16 */
                {8'hee,8'hxx} : dec_pc_inc3 = 1'b1;  /* BR,,$!addr16 */
                {8'h61,8'hc3} : dec_pc_inc3 = 1'b1;  /* BH,,$addr8 */
                {8'h61,8'hd3} : dec_pc_inc3 = 1'b1;  /* BNH,,$addr8 */
                {8'h31,8'h03} : dec_pc_inc3 = 1'b1;  /* BT,A.0,$addr8 */
                {8'h31,8'h13} : dec_pc_inc3 = 1'b1;  /* BT,A.1,$addr8 */
                {8'h31,8'h23} : dec_pc_inc3 = 1'b1;  /* BT,A.2,$addr8 */
                {8'h31,8'h33} : dec_pc_inc3 = 1'b1;  /* BT,A.3,$addr8 */
                {8'h31,8'h43} : dec_pc_inc3 = 1'b1;  /* BT,A.4,$addr8 */
                {8'h31,8'h53} : dec_pc_inc3 = 1'b1;  /* BT,A.5,$addr8 */
                {8'h31,8'h63} : dec_pc_inc3 = 1'b1;  /* BT,A.6,$addr8 */
                {8'h31,8'h73} : dec_pc_inc3 = 1'b1;  /* BT,A.7,$addr8 */
                {8'h31,8'h83} : dec_pc_inc3 = 1'b1;  /* BT,[HL].0,$addr8 */
                {8'h31,8'h93} : dec_pc_inc3 = 1'b1;  /* BT,[HL].1,$addr8 */
                {8'h31,8'ha3} : dec_pc_inc3 = 1'b1;  /* BT,[HL].2,$addr8 */
                {8'h31,8'hb3} : dec_pc_inc3 = 1'b1;  /* BT,[HL].3,$addr8 */
                {8'h31,8'hc3} : dec_pc_inc3 = 1'b1;  /* BT,[HL].4,$addr8 */
                {8'h31,8'hd3} : dec_pc_inc3 = 1'b1;  /* BT,[HL].5,$addr8 */
                {8'h31,8'he3} : dec_pc_inc3 = 1'b1;  /* BT,[HL].6,$addr8 */
                {8'h31,8'hf3} : dec_pc_inc3 = 1'b1;  /* BT,[HL].7,$addr8 */
                {8'h31,8'h05} : dec_pc_inc3 = 1'b1;  /* BF,A.0,$addr8 */
                {8'h31,8'h15} : dec_pc_inc3 = 1'b1;  /* BF,A.1,$addr8 */
                {8'h31,8'h25} : dec_pc_inc3 = 1'b1;  /* BF,A.2,$addr8 */
                {8'h31,8'h35} : dec_pc_inc3 = 1'b1;  /* BF,A.3,$addr8 */
                {8'h31,8'h45} : dec_pc_inc3 = 1'b1;  /* BF,A.4,$addr8 */
                {8'h31,8'h55} : dec_pc_inc3 = 1'b1;  /* BF,A.5,$addr8 */
                {8'h31,8'h65} : dec_pc_inc3 = 1'b1;  /* BF,A.6,$addr8 */
                {8'h31,8'h75} : dec_pc_inc3 = 1'b1;  /* BF,A.7,$addr8 */
                {8'h31,8'h85} : dec_pc_inc3 = 1'b1;  /* BF,[HL].0,$addr8 */
                {8'h31,8'h95} : dec_pc_inc3 = 1'b1;  /* BF,[HL].1,$addr8 */
                {8'h31,8'ha5} : dec_pc_inc3 = 1'b1;  /* BF,[HL].2,$addr8 */
                {8'h31,8'hb5} : dec_pc_inc3 = 1'b1;  /* BF,[HL].3,$addr8 */
                {8'h31,8'hc5} : dec_pc_inc3 = 1'b1;  /* BF,[HL].4,$addr8 */
                {8'h31,8'hd5} : dec_pc_inc3 = 1'b1;  /* BF,[HL].5,$addr8 */
                {8'h31,8'he5} : dec_pc_inc3 = 1'b1;  /* BF,[HL].6,$addr8 */
                {8'h31,8'hf5} : dec_pc_inc3 = 1'b1;  /* BF,[HL].7,$addr8 */
                {8'h31,8'h01} : dec_pc_inc3 = 1'b1;  /* BTCLR,A.0,$addr8 */
                {8'h31,8'h11} : dec_pc_inc3 = 1'b1;  /* BTCLR,A.1,$addr8 */
                {8'h31,8'h21} : dec_pc_inc3 = 1'b1;  /* BTCLR,A.2,$addr8 */
                {8'h31,8'h31} : dec_pc_inc3 = 1'b1;  /* BTCLR,A.3,$addr8 */
                {8'h31,8'h41} : dec_pc_inc3 = 1'b1;  /* BTCLR,A.4,$addr8 */
                {8'h31,8'h51} : dec_pc_inc3 = 1'b1;  /* BTCLR,A.5,$addr8 */
                {8'h31,8'h61} : dec_pc_inc3 = 1'b1;  /* BTCLR,A.6,$addr8 */
                {8'h31,8'h71} : dec_pc_inc3 = 1'b1;  /* BTCLR,A.7,$addr8 */
                {8'h31,8'h81} : dec_pc_inc3 = 1'b1;  /* BTCLR,[HL].0,$addr8 */
                {8'h31,8'h91} : dec_pc_inc3 = 1'b1;  /* BTCLR,[HL].1,$addr8 */
                {8'h31,8'ha1} : dec_pc_inc3 = 1'b1;  /* BTCLR,[HL].2,$addr8 */
                {8'h31,8'hb1} : dec_pc_inc3 = 1'b1;  /* BTCLR,[HL].3,$addr8 */
                {8'h31,8'hc1} : dec_pc_inc3 = 1'b1;  /* BTCLR,[HL].4,$addr8 */
                {8'h31,8'hd1} : dec_pc_inc3 = 1'b1;  /* BTCLR,[HL].5,$addr8 */
                {8'h31,8'he1} : dec_pc_inc3 = 1'b1;  /* BTCLR,[HL].6,$addr8 */
                {8'h31,8'hf1} : dec_pc_inc3 = 1'b1;  /* BTCLR,[HL].7,$addr8 */
                {8'h61,8'hb1} : dec_pc_inc3 = 1'b1;  /* SOFT3,,BREAK */
                {8'h61,8'hbb} : dec_pc_inc3 = 1'b1;  /* XCH,A,sfr */
                {8'h61,8'hbf} : dec_pc_inc3 = 1'b1;  /* XCH,A,[DE+byte] */
                {8'h61,8'hbd} : dec_pc_inc3 = 1'b1;  /* XCH,A,[HL+byte] */
                default : dec_pc_inc3 = 1'b0;
            endcase
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'hcd,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV,saddr,#byte */
                {8'hce,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV,sfr,#byte */
                {8'hca,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV,[DE+byte],#byte */
                {8'hcc,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV,[HL+byte],#byte */
                {8'h8f,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV,A,!addr16 */
                {8'h9f,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV,!addr16,A */
                {8'h09,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV,A,word[B] */
                {8'h18,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV,word[B],A */
                {8'h29,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV,A,word[C] */
                {8'h28,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV,word[C],A */
                {8'h49,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV,A,word[BC] */
                {8'h48,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV,word[BC],A */
                {8'hc8,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV,[SP+byte],#byte */
                {8'he9,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV,B,!addr16 */
                {8'hf9,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV,C,!addr16 */
                {8'hd9,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV,X,!addr16 */
                {8'h61,8'hb8,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV,ES,saddr */
                {8'h61,8'hce,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOVS,[HL+byte],X */
                {8'h61,8'ha8,2'bx1} : dec_pc_inc3 = 1'b1;  /* XCH,A,saddr */
                {8'h61,8'hab,2'bx1} : dec_pc_inc3 = 1'b1;  /* XCH,A,sfr */
                {8'h61,8'haf,2'bx1} : dec_pc_inc3 = 1'b1;  /* XCH,A,[DE+byte] */
                {8'h61,8'had,2'bx1} : dec_pc_inc3 = 1'b1;  /* XCH,A,[HL+byte] */
                {8'he5,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* ONEB,,!addr16 */
                {8'hf5,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* CLRB,,!addr16 */
                {8'h30,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOVW,AX,#word */
                {8'h32,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOVW,BC,#word */
                {8'h34,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOVW,DE,#word */
                {8'h36,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOVW,HL,#word */
                {8'haf,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOVW,AX,!addr16 */
                {8'hbf,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOVW,!addr16,AX */
                {8'h59,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOVW,AX,word[B] */
                {8'h58,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOVW,word[B],AX */
                {8'h69,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOVW,AX,word[C] */
                {8'h68,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOVW,word[C],AX */
                {8'h79,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOVW,AX,word[BC] */
                {8'h78,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOVW,word[BC],AX */
                {8'hdb,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOVW,BC,!addr16 */
                {8'heb,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOVW,DE,!addr16 */
                {8'hfb,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOVW,HL,!addr16 */
                {8'h0a,8'hxx,2'bx1} : dec_pc_inc3 = 1'b1;  /* ADD,saddr,#byte */
                {8'h0f,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* ADD,A,!addr16 */
                {8'h1a,8'hxx,2'bx1} : dec_pc_inc3 = 1'b1;  /* ADDC,saddr,#byte */
                {8'h1f,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* ADDC,A,!addr16 */
                {8'h2a,8'hxx,2'bx1} : dec_pc_inc3 = 1'b1;  /* SUB,saddr,#byte */
                {8'h2f,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* SUB,A,!addr16 */
                {8'h3a,8'hxx,2'bx1} : dec_pc_inc3 = 1'b1;  /* SUBC,saddr,#byte */
                {8'h3f,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* SUBC,A,!addr16 */
                {8'h5a,8'hxx,2'bx1} : dec_pc_inc3 = 1'b1;  /* AND,saddr,#byte */
                {8'h5f,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* AND,A,!addr16 */
                {8'h6a,8'hxx,2'bx1} : dec_pc_inc3 = 1'b1;  /* OR,saddr,#byte */
                {8'h6f,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* OR,A,!addr16 */
                {8'h7a,8'hxx,2'bx1} : dec_pc_inc3 = 1'b1;  /* XOR,saddr,#byte */
                {8'h7f,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* XOR,A,!addr16 */
                {8'h4a,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* CMP,saddr,#byte */
                {8'h4f,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* CMP,A,!addr16 */
                {8'h61,8'hde,2'bxx} : dec_pc_inc3 = 1'b1;  /* CMPS,X,[HL+byte] */
                {8'hd5,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* CMP0,,!addr16 */
                {8'h04,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* ADDW,AX,#word */
                {8'h02,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* ADDW,AX,!addr16 */
                {8'h61,8'h09,2'bxx} : dec_pc_inc3 = 1'b1;  /* ADDW,AX,[HL+byte] */
                {8'h24,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* SUBW,AX,#word */
                {8'h22,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* SUBW,AX,!addr16 */
                {8'h61,8'h29,2'bxx} : dec_pc_inc3 = 1'b1;  /* SUBW,AX,[HL+byte] */
                {8'h44,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* CMPW,AX,#word */
                {8'h42,8'hxx,2'bxx} : dec_pc_inc3 = 1'b1;  /* CMPW,AX,!addr16 */
                {8'h61,8'h49,2'bxx} : dec_pc_inc3 = 1'b1;  /* CMPW,AX,[HL+byte] */
                {8'ha0,8'hxx,2'bx1} : dec_pc_inc3 = 1'b1;  /* INC,,!addr16 */
                {8'h61,8'h59,2'bx1} : dec_pc_inc3 = 1'b1;  /* INC,,[HL+byte] */
                {8'hb0,8'hxx,2'bx1} : dec_pc_inc3 = 1'b1;  /* DEC,,!addr16 */
                {8'h61,8'h69,2'bx1} : dec_pc_inc3 = 1'b1;  /* DEC,,[HL+byte] */
                {8'ha2,8'hxx,2'bx1} : dec_pc_inc3 = 1'b1;  /* INCW,,!addr16 */
                {8'h61,8'h79,2'bx1} : dec_pc_inc3 = 1'b1;  /* INCW,,[HL+byte] */
                {8'hb2,8'hxx,2'bx1} : dec_pc_inc3 = 1'b1;  /* DECW,,!addr16 */
                {8'h61,8'h89,2'bx1} : dec_pc_inc3 = 1'b1;  /* DECW,,[HL+byte] */
                {8'h71,8'h04,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,saddr.0 */
                {8'h71,8'h14,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,saddr.1 */
                {8'h71,8'h24,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,saddr.2 */
                {8'h71,8'h34,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,saddr.3 */
                {8'h71,8'h44,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,saddr.4 */
                {8'h71,8'h54,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,saddr.5 */
                {8'h71,8'h64,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,saddr.6 */
                {8'h71,8'h74,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,saddr.7 */
                {8'h71,8'h0c,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,sfr.0 */
                {8'h71,8'h1c,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,sfr.1 */
                {8'h71,8'h2c,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,sfr.2 */
                {8'h71,8'h3c,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,sfr.3 */
                {8'h71,8'h4c,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,sfr.4 */
                {8'h71,8'h5c,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,sfr.5 */
                {8'h71,8'h6c,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,sfr.6 */
                {8'h71,8'h7c,2'bxx} : dec_pc_inc3 = 1'b1;  /* MOV1,CY,sfr.7 */
                {8'h71,8'h01,2'bx1} : dec_pc_inc3 = 1'b1;  /* MOV1,saddr.0,CY */
                {8'h71,8'h11,2'bx1} : dec_pc_inc3 = 1'b1;  /* MOV1,saddr.1,CY */
                {8'h71,8'h21,2'bx1} : dec_pc_inc3 = 1'b1;  /* MOV1,saddr.2,CY */
                {8'h71,8'h31,2'bx1} : dec_pc_inc3 = 1'b1;  /* MOV1,saddr.3,CY */
                {8'h71,8'h41,2'bx1} : dec_pc_inc3 = 1'b1;  /* MOV1,saddr.4,CY */
                {8'h71,8'h51,2'bx1} : dec_pc_inc3 = 1'b1;  /* MOV1,saddr.5,CY */
                {8'h71,8'h61,2'bx1} : dec_pc_inc3 = 1'b1;  /* MOV1,saddr.6,CY */
                {8'h71,8'h71,2'bx1} : dec_pc_inc3 = 1'b1;  /* MOV1,saddr.7,CY */
                {8'h71,8'h09,2'bx1} : dec_pc_inc3 = 1'b1;  /* MOV1,sfr.0,CY */
                {8'h71,8'h19,2'bx1} : dec_pc_inc3 = 1'b1;  /* MOV1,sfr.1,CY */
                {8'h71,8'h29,2'bx1} : dec_pc_inc3 = 1'b1;  /* MOV1,sfr.2,CY */
                {8'h71,8'h39,2'bx1} : dec_pc_inc3 = 1'b1;  /* MOV1,sfr.3,CY */
                {8'h71,8'h49,2'bx1} : dec_pc_inc3 = 1'b1;  /* MOV1,sfr.4,CY */
                {8'h71,8'h59,2'bx1} : dec_pc_inc3 = 1'b1;  /* MOV1,sfr.5,CY */
                {8'h71,8'h69,2'bx1} : dec_pc_inc3 = 1'b1;  /* MOV1,sfr.6,CY */
                {8'h71,8'h79,2'bx1} : dec_pc_inc3 = 1'b1;  /* MOV1,sfr.7,CY */
                {8'h71,8'h05,2'bxx} : dec_pc_inc3 = 1'b1;  /* AND1,CY,saddr.0 */
                {8'h71,8'h15,2'bxx} : dec_pc_inc3 = 1'b1;  /* AND1,CY,saddr.1 */
                {8'h71,8'h25,2'bxx} : dec_pc_inc3 = 1'b1;  /* AND1,CY,saddr.2 */
                {8'h71,8'h35,2'bxx} : dec_pc_inc3 = 1'b1;  /* AND1,CY,saddr.3 */
                {8'h71,8'h45,2'bxx} : dec_pc_inc3 = 1'b1;  /* AND1,CY,saddr.4 */
                {8'h71,8'h55,2'bxx} : dec_pc_inc3 = 1'b1;  /* AND1,CY,saddr.5 */
                {8'h71,8'h65,2'bxx} : dec_pc_inc3 = 1'b1;  /* AND1,CY,saddr.6 */
                {8'h71,8'h75,2'bxx} : dec_pc_inc3 = 1'b1;  /* AND1,CY,saddr.7 */
                {8'h71,8'h0d,2'bxx} : dec_pc_inc3 = 1'b1;  /* AND1,CY,sfr.0 */
                {8'h71,8'h1d,2'bxx} : dec_pc_inc3 = 1'b1;  /* AND1,CY,sfr.1 */
                {8'h71,8'h2d,2'bxx} : dec_pc_inc3 = 1'b1;  /* AND1,CY,sfr.2 */
                {8'h71,8'h3d,2'bxx} : dec_pc_inc3 = 1'b1;  /* AND1,CY,sfr.3 */
                {8'h71,8'h4d,2'bxx} : dec_pc_inc3 = 1'b1;  /* AND1,CY,sfr.4 */
                {8'h71,8'h5d,2'bxx} : dec_pc_inc3 = 1'b1;  /* AND1,CY,sfr.5 */
                {8'h71,8'h6d,2'bxx} : dec_pc_inc3 = 1'b1;  /* AND1,CY,sfr.6 */
                {8'h71,8'h7d,2'bxx} : dec_pc_inc3 = 1'b1;  /* AND1,CY,sfr.7 */
                {8'h71,8'h06,2'bxx} : dec_pc_inc3 = 1'b1;  /* OR1,CY,saddr.0 */
                {8'h71,8'h16,2'bxx} : dec_pc_inc3 = 1'b1;  /* OR1,CY,saddr.1 */
                {8'h71,8'h26,2'bxx} : dec_pc_inc3 = 1'b1;  /* OR1,CY,saddr.2 */
                {8'h71,8'h36,2'bxx} : dec_pc_inc3 = 1'b1;  /* OR1,CY,saddr.3 */
                {8'h71,8'h46,2'bxx} : dec_pc_inc3 = 1'b1;  /* OR1,CY,saddr.4 */
                {8'h71,8'h56,2'bxx} : dec_pc_inc3 = 1'b1;  /* OR1,CY,saddr.5 */
                {8'h71,8'h66,2'bxx} : dec_pc_inc3 = 1'b1;  /* OR1,CY,saddr.6 */
                {8'h71,8'h76,2'bxx} : dec_pc_inc3 = 1'b1;  /* OR1,CY,saddr.7 */
                {8'h71,8'h0e,2'bxx} : dec_pc_inc3 = 1'b1;  /* OR1,CY,sfr.0 */
                {8'h71,8'h1e,2'bxx} : dec_pc_inc3 = 1'b1;  /* OR1,CY,sfr.1 */
                {8'h71,8'h2e,2'bxx} : dec_pc_inc3 = 1'b1;  /* OR1,CY,sfr.2 */
                {8'h71,8'h3e,2'bxx} : dec_pc_inc3 = 1'b1;  /* OR1,CY,sfr.3 */
                {8'h71,8'h4e,2'bxx} : dec_pc_inc3 = 1'b1;  /* OR1,CY,sfr.4 */
                {8'h71,8'h5e,2'bxx} : dec_pc_inc3 = 1'b1;  /* OR1,CY,sfr.5 */
                {8'h71,8'h6e,2'bxx} : dec_pc_inc3 = 1'b1;  /* OR1,CY,sfr.6 */
                {8'h71,8'h7e,2'bxx} : dec_pc_inc3 = 1'b1;  /* OR1,CY,sfr.7 */
                {8'h71,8'h07,2'bxx} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,saddr.0 */
                {8'h71,8'h17,2'bxx} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,saddr.1 */
                {8'h71,8'h27,2'bxx} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,saddr.2 */
                {8'h71,8'h37,2'bxx} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,saddr.3 */
                {8'h71,8'h47,2'bxx} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,saddr.4 */
                {8'h71,8'h57,2'bxx} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,saddr.5 */
                {8'h71,8'h67,2'bxx} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,saddr.6 */
                {8'h71,8'h77,2'bxx} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,saddr.7 */
                {8'h71,8'h0f,2'bxx} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,sfr.0 */
                {8'h71,8'h1f,2'bxx} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,sfr.1 */
                {8'h71,8'h2f,2'bxx} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,sfr.2 */
                {8'h71,8'h3f,2'bxx} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,sfr.3 */
                {8'h71,8'h4f,2'bxx} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,sfr.4 */
                {8'h71,8'h5f,2'bxx} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,sfr.5 */
                {8'h71,8'h6f,2'bxx} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,sfr.6 */
                {8'h71,8'h7f,2'bxx} : dec_pc_inc3 = 1'b1;  /* XOR1,CY,sfr.7 */
                {8'h71,8'h02,2'bx1} : dec_pc_inc3 = 1'b1;  /* SET1,,saddr.0 */
                {8'h71,8'h12,2'bx1} : dec_pc_inc3 = 1'b1;  /* SET1,,saddr.1 */
                {8'h71,8'h22,2'bx1} : dec_pc_inc3 = 1'b1;  /* SET1,,saddr.2 */
                {8'h71,8'h32,2'bx1} : dec_pc_inc3 = 1'b1;  /* SET1,,saddr.3 */
                {8'h71,8'h42,2'bx1} : dec_pc_inc3 = 1'b1;  /* SET1,,saddr.4 */
                {8'h71,8'h52,2'bx1} : dec_pc_inc3 = 1'b1;  /* SET1,,saddr.5 */
                {8'h71,8'h62,2'bx1} : dec_pc_inc3 = 1'b1;  /* SET1,,saddr.6 */
                {8'h71,8'h72,2'bx1} : dec_pc_inc3 = 1'b1;  /* SET1,,saddr.7 */
                {8'h71,8'h0a,2'bx1} : dec_pc_inc3 = 1'b1;  /* SET1,,sfr.0 */
                {8'h71,8'h1a,2'bx1} : dec_pc_inc3 = 1'b1;  /* SET1,,sfr.1 */
                {8'h71,8'h2a,2'bx1} : dec_pc_inc3 = 1'b1;  /* SET1,,sfr.2 */
                {8'h71,8'h3a,2'bx1} : dec_pc_inc3 = 1'b1;  /* SET1,,sfr.3 */
                {8'h71,8'h4a,2'bx1} : dec_pc_inc3 = 1'b1;  /* SET1,,sfr.4 */
                {8'h71,8'h5a,2'bx1} : dec_pc_inc3 = 1'b1;  /* SET1,,sfr.5 */
                {8'h71,8'h6a,2'bx1} : dec_pc_inc3 = 1'b1;  /* SET1,,sfr.6 */
                {8'h71,8'h7a,2'bx1} : dec_pc_inc3 = 1'b1;  /* SET1,,sfr.7 */
                {8'h71,8'h03,2'bx1} : dec_pc_inc3 = 1'b1;  /* CLR1,,saddr.0 */
                {8'h71,8'h13,2'bx1} : dec_pc_inc3 = 1'b1;  /* CLR1,,saddr.1 */
                {8'h71,8'h23,2'bx1} : dec_pc_inc3 = 1'b1;  /* CLR1,,saddr.2 */
                {8'h71,8'h33,2'bx1} : dec_pc_inc3 = 1'b1;  /* CLR1,,saddr.3 */
                {8'h71,8'h43,2'bx1} : dec_pc_inc3 = 1'b1;  /* CLR1,,saddr.4 */
                {8'h71,8'h53,2'bx1} : dec_pc_inc3 = 1'b1;  /* CLR1,,saddr.5 */
                {8'h71,8'h63,2'bx1} : dec_pc_inc3 = 1'b1;  /* CLR1,,saddr.6 */
                {8'h71,8'h73,2'bx1} : dec_pc_inc3 = 1'b1;  /* CLR1,,saddr.7 */
                {8'h71,8'h0b,2'bx1} : dec_pc_inc3 = 1'b1;  /* CLR1,,sfr.0 */
                {8'h71,8'h1b,2'bx1} : dec_pc_inc3 = 1'b1;  /* CLR1,,sfr.1 */
                {8'h71,8'h2b,2'bx1} : dec_pc_inc3 = 1'b1;  /* CLR1,,sfr.2 */
                {8'h71,8'h3b,2'bx1} : dec_pc_inc3 = 1'b1;  /* CLR1,,sfr.3 */
                {8'h71,8'h4b,2'bx1} : dec_pc_inc3 = 1'b1;  /* CLR1,,sfr.4 */
                {8'h71,8'h5b,2'bx1} : dec_pc_inc3 = 1'b1;  /* CLR1,,sfr.5 */
                {8'h71,8'h6b,2'bx1} : dec_pc_inc3 = 1'b1;  /* CLR1,,sfr.6 */
                {8'h71,8'h7b,2'bx1} : dec_pc_inc3 = 1'b1;  /* CLR1,,sfr.7 */
                {8'hfe,8'hxx,2'bx0} : dec_pc_inc3 = 1'b1;  /* CALL,,$!addr16 */
                {8'hfd,8'hxx,2'bx0} : dec_pc_inc3 = 1'b1;  /* CALL,,!addr16 */
                {8'hee,8'hxx,2'bx0} : dec_pc_inc3 = 1'b1;  /* BR,,$!addr16 */
                {8'h61,8'hc3,2'bx1} : dec_pc_inc3 = 1'b1;  /* BH,,$addr8 */
                {8'h61,8'hd3,2'bx1} : dec_pc_inc3 = 1'b1;  /* BNH,,$addr8 */
                {8'h31,8'h03,2'b10} : dec_pc_inc3 = 1'b1;  /* BT,A.0,$addr8 */
                {8'h31,8'h13,2'b10} : dec_pc_inc3 = 1'b1;  /* BT,A.1,$addr8 */
                {8'h31,8'h23,2'b10} : dec_pc_inc3 = 1'b1;  /* BT,A.2,$addr8 */
                {8'h31,8'h33,2'b10} : dec_pc_inc3 = 1'b1;  /* BT,A.3,$addr8 */
                {8'h31,8'h43,2'b10} : dec_pc_inc3 = 1'b1;  /* BT,A.4,$addr8 */
                {8'h31,8'h53,2'b10} : dec_pc_inc3 = 1'b1;  /* BT,A.5,$addr8 */
                {8'h31,8'h63,2'b10} : dec_pc_inc3 = 1'b1;  /* BT,A.6,$addr8 */
                {8'h31,8'h73,2'b10} : dec_pc_inc3 = 1'b1;  /* BT,A.7,$addr8 */
                {8'h31,8'h83,2'b10} : dec_pc_inc3 = 1'b1;  /* BT,[HL].0,$addr8 */
                {8'h31,8'h93,2'b10} : dec_pc_inc3 = 1'b1;  /* BT,[HL].1,$addr8 */
                {8'h31,8'ha3,2'b10} : dec_pc_inc3 = 1'b1;  /* BT,[HL].2,$addr8 */
                {8'h31,8'hb3,2'b10} : dec_pc_inc3 = 1'b1;  /* BT,[HL].3,$addr8 */
                {8'h31,8'hc3,2'b10} : dec_pc_inc3 = 1'b1;  /* BT,[HL].4,$addr8 */
                {8'h31,8'hd3,2'b10} : dec_pc_inc3 = 1'b1;  /* BT,[HL].5,$addr8 */
                {8'h31,8'he3,2'b10} : dec_pc_inc3 = 1'b1;  /* BT,[HL].6,$addr8 */
                {8'h31,8'hf3,2'b10} : dec_pc_inc3 = 1'b1;  /* BT,[HL].7,$addr8 */
                {8'h31,8'h05,2'b10} : dec_pc_inc3 = 1'b1;  /* BF,A.0,$addr8 */
                {8'h31,8'h15,2'b10} : dec_pc_inc3 = 1'b1;  /* BF,A.1,$addr8 */
                {8'h31,8'h25,2'b10} : dec_pc_inc3 = 1'b1;  /* BF,A.2,$addr8 */
                {8'h31,8'h35,2'b10} : dec_pc_inc3 = 1'b1;  /* BF,A.3,$addr8 */
                {8'h31,8'h45,2'b10} : dec_pc_inc3 = 1'b1;  /* BF,A.4,$addr8 */
                {8'h31,8'h55,2'b10} : dec_pc_inc3 = 1'b1;  /* BF,A.5,$addr8 */
                {8'h31,8'h65,2'b10} : dec_pc_inc3 = 1'b1;  /* BF,A.6,$addr8 */
                {8'h31,8'h75,2'b10} : dec_pc_inc3 = 1'b1;  /* BF,A.7,$addr8 */
                {8'h31,8'h85,2'b10} : dec_pc_inc3 = 1'b1;  /* BF,[HL].0,$addr8 */
                {8'h31,8'h95,2'b10} : dec_pc_inc3 = 1'b1;  /* BF,[HL].1,$addr8 */
                {8'h31,8'ha5,2'b10} : dec_pc_inc3 = 1'b1;  /* BF,[HL].2,$addr8 */
                {8'h31,8'hb5,2'b10} : dec_pc_inc3 = 1'b1;  /* BF,[HL].3,$addr8 */
                {8'h31,8'hc5,2'b10} : dec_pc_inc3 = 1'b1;  /* BF,[HL].4,$addr8 */
                {8'h31,8'hd5,2'b10} : dec_pc_inc3 = 1'b1;  /* BF,[HL].5,$addr8 */
                {8'h31,8'he5,2'b10} : dec_pc_inc3 = 1'b1;  /* BF,[HL].6,$addr8 */
                {8'h31,8'hf5,2'b10} : dec_pc_inc3 = 1'b1;  /* BF,[HL].7,$addr8 */
                {8'h31,8'h01,2'b10} : dec_pc_inc3 = 1'b1;  /* BTCLR,A.0,$addr8 */
                {8'h31,8'h11,2'b10} : dec_pc_inc3 = 1'b1;  /* BTCLR,A.1,$addr8 */
                {8'h31,8'h21,2'b10} : dec_pc_inc3 = 1'b1;  /* BTCLR,A.2,$addr8 */
                {8'h31,8'h31,2'b10} : dec_pc_inc3 = 1'b1;  /* BTCLR,A.3,$addr8 */
                {8'h31,8'h41,2'b10} : dec_pc_inc3 = 1'b1;  /* BTCLR,A.4,$addr8 */
                {8'h31,8'h51,2'b10} : dec_pc_inc3 = 1'b1;  /* BTCLR,A.5,$addr8 */
                {8'h31,8'h61,2'b10} : dec_pc_inc3 = 1'b1;  /* BTCLR,A.6,$addr8 */
                {8'h31,8'h71,2'b10} : dec_pc_inc3 = 1'b1;  /* BTCLR,A.7,$addr8 */
                {8'h31,8'h81,2'b10} : dec_pc_inc3 = 1'b1;  /* BTCLR,[HL].0,$addr8 */
                {8'h31,8'h91,2'b10} : dec_pc_inc3 = 1'b1;  /* BTCLR,[HL].1,$addr8 */
                {8'h31,8'ha1,2'b10} : dec_pc_inc3 = 1'b1;  /* BTCLR,[HL].2,$addr8 */
                {8'h31,8'hb1,2'b10} : dec_pc_inc3 = 1'b1;  /* BTCLR,[HL].3,$addr8 */
                {8'h31,8'hc1,2'b10} : dec_pc_inc3 = 1'b1;  /* BTCLR,[HL].4,$addr8 */
                {8'h31,8'hd1,2'b10} : dec_pc_inc3 = 1'b1;  /* BTCLR,[HL].5,$addr8 */
                {8'h31,8'he1,2'b10} : dec_pc_inc3 = 1'b1;  /* BTCLR,[HL].6,$addr8 */
                {8'h31,8'hf1,2'b10} : dec_pc_inc3 = 1'b1;  /* BTCLR,[HL].7,$addr8 */
                {8'h61,8'hb1,2'bx0} : dec_pc_inc3 = 1'b1;  /* SOFT3,,BREAK */
                {8'h61,8'hbb,2'bx1} : dec_pc_inc3 = 1'b1;  /* XCH,A,sfr */
                {8'h61,8'hbf,2'bx1} : dec_pc_inc3 = 1'b1;  /* XCH,A,[DE+byte] */
                {8'h61,8'hbd,2'bx1} : dec_pc_inc3 = 1'b1;  /* XCH,A,[HL+byte] */
                default : dec_pc_inc3 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_pc_inc4;
    reg    dec_pc_inc4;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1) begin
            dec_pc_inc4 = 1'b0;
        end else if(skpack == 1'b1) begin
            casex ({ID_stage0,ID_stage1})  
                {8'hcf,8'hxx} : dec_pc_inc4 = 1'b1;  /* MOV,!addr16,#byte */
                {8'h19,8'hxx} : dec_pc_inc4 = 1'b1;  /* MOV,word[B],#byte */
                {8'h38,8'hxx} : dec_pc_inc4 = 1'b1;  /* MOV,word[C],#byte */
                {8'h39,8'hxx} : dec_pc_inc4 = 1'b1;  /* MOV,word[BC],#byte */
                {8'h61,8'haa} : dec_pc_inc4 = 1'b1;  /* XCH,A,!addr16 */
                {8'hc9,8'hxx} : dec_pc_inc4 = 1'b1;  /* MOVW,saddrp,#word */
                {8'hcb,8'hxx} : dec_pc_inc4 = 1'b1;  /* MOVW,sfrp,#word */
                {8'h40,8'hxx} : dec_pc_inc4 = 1'b1;  /* CMP,!addr16,#byte */
                {8'h71,8'h00} : dec_pc_inc4 = 1'b1;  /* SET1,,!addr16.0 */
                {8'h71,8'h10} : dec_pc_inc4 = 1'b1;  /* SET1,,!addr16.1 */
                {8'h71,8'h20} : dec_pc_inc4 = 1'b1;  /* SET1,,!addr16.2 */
                {8'h71,8'h30} : dec_pc_inc4 = 1'b1;  /* SET1,,!addr16.3 */
                {8'h71,8'h40} : dec_pc_inc4 = 1'b1;  /* SET1,,!addr16.4 */
                {8'h71,8'h50} : dec_pc_inc4 = 1'b1;  /* SET1,,!addr16.5 */
                {8'h71,8'h60} : dec_pc_inc4 = 1'b1;  /* SET1,,!addr16.6 */
                {8'h71,8'h70} : dec_pc_inc4 = 1'b1;  /* SET1,,!addr16.7 */
                {8'h71,8'h08} : dec_pc_inc4 = 1'b1;  /* CLR1,,!addr16.0 */
                {8'h71,8'h18} : dec_pc_inc4 = 1'b1;  /* CLR1,,!addr16.1 */
                {8'h71,8'h28} : dec_pc_inc4 = 1'b1;  /* CLR1,,!addr16.2 */
                {8'h71,8'h38} : dec_pc_inc4 = 1'b1;  /* CLR1,,!addr16.3 */
                {8'h71,8'h48} : dec_pc_inc4 = 1'b1;  /* CLR1,,!addr16.4 */
                {8'h71,8'h58} : dec_pc_inc4 = 1'b1;  /* CLR1,,!addr16.5 */
                {8'h71,8'h68} : dec_pc_inc4 = 1'b1;  /* CLR1,,!addr16.6 */
                {8'h71,8'h78} : dec_pc_inc4 = 1'b1;  /* CLR1,,!addr16.7 */
                {8'hfc,8'hxx} : dec_pc_inc4 = 1'b1;  /* CALL,,!!addr20 */
                {8'hec,8'hxx} : dec_pc_inc4 = 1'b1;  /* BR,,!!addr20 */
                {8'h31,8'h02} : dec_pc_inc4 = 1'b1;  /* BT,saddr.0,$addr8 */
                {8'h31,8'h12} : dec_pc_inc4 = 1'b1;  /* BT,saddr.1,$addr8 */
                {8'h31,8'h22} : dec_pc_inc4 = 1'b1;  /* BT,saddr.2,$addr8 */
                {8'h31,8'h32} : dec_pc_inc4 = 1'b1;  /* BT,saddr.3,$addr8 */
                {8'h31,8'h42} : dec_pc_inc4 = 1'b1;  /* BT,saddr.4,$addr8 */
                {8'h31,8'h52} : dec_pc_inc4 = 1'b1;  /* BT,saddr.5,$addr8 */
                {8'h31,8'h62} : dec_pc_inc4 = 1'b1;  /* BT,saddr.6,$addr8 */
                {8'h31,8'h72} : dec_pc_inc4 = 1'b1;  /* BT,saddr.7,$addr8 */
                {8'h31,8'h82} : dec_pc_inc4 = 1'b1;  /* BT,sfr.0,$addr8 */
                {8'h31,8'h92} : dec_pc_inc4 = 1'b1;  /* BT,sfr.1,$addr8 */
                {8'h31,8'ha2} : dec_pc_inc4 = 1'b1;  /* BT,sfr.2,$addr8 */
                {8'h31,8'hb2} : dec_pc_inc4 = 1'b1;  /* BT,sfr.3,$addr8 */
                {8'h31,8'hc2} : dec_pc_inc4 = 1'b1;  /* BT,sfr.4,$addr8 */
                {8'h31,8'hd2} : dec_pc_inc4 = 1'b1;  /* BT,sfr.5,$addr8 */
                {8'h31,8'he2} : dec_pc_inc4 = 1'b1;  /* BT,sfr.6,$addr8 */
                {8'h31,8'hf2} : dec_pc_inc4 = 1'b1;  /* BT,sfr.7,$addr8 */
                {8'h31,8'h04} : dec_pc_inc4 = 1'b1;  /* BF,saddr.0,$addr8 */
                {8'h31,8'h14} : dec_pc_inc4 = 1'b1;  /* BF,saddr.1,$addr8 */
                {8'h31,8'h24} : dec_pc_inc4 = 1'b1;  /* BF,saddr.2,$addr8 */
                {8'h31,8'h34} : dec_pc_inc4 = 1'b1;  /* BF,saddr.3,$addr8 */
                {8'h31,8'h44} : dec_pc_inc4 = 1'b1;  /* BF,saddr.4,$addr8 */
                {8'h31,8'h54} : dec_pc_inc4 = 1'b1;  /* BF,saddr.5,$addr8 */
                {8'h31,8'h64} : dec_pc_inc4 = 1'b1;  /* BF,saddr.6,$addr8 */
                {8'h31,8'h74} : dec_pc_inc4 = 1'b1;  /* BF,saddr.7,$addr8 */
                {8'h31,8'h84} : dec_pc_inc4 = 1'b1;  /* BF,sfr.0,$addr8 */
                {8'h31,8'h94} : dec_pc_inc4 = 1'b1;  /* BF,sfr.1,$addr8 */
                {8'h31,8'ha4} : dec_pc_inc4 = 1'b1;  /* BF,sfr.2,$addr8 */
                {8'h31,8'hb4} : dec_pc_inc4 = 1'b1;  /* BF,sfr.3,$addr8 */
                {8'h31,8'hc4} : dec_pc_inc4 = 1'b1;  /* BF,sfr.4,$addr8 */
                {8'h31,8'hd4} : dec_pc_inc4 = 1'b1;  /* BF,sfr.5,$addr8 */
                {8'h31,8'he4} : dec_pc_inc4 = 1'b1;  /* BF,sfr.6,$addr8 */
                {8'h31,8'hf4} : dec_pc_inc4 = 1'b1;  /* BF,sfr.7,$addr8 */
                {8'h31,8'h00} : dec_pc_inc4 = 1'b1;  /* BTCLR,saddr.0,$addr8 */
                {8'h31,8'h10} : dec_pc_inc4 = 1'b1;  /* BTCLR,saddr.1,$addr8 */
                {8'h31,8'h20} : dec_pc_inc4 = 1'b1;  /* BTCLR,saddr.2,$addr8 */
                {8'h31,8'h30} : dec_pc_inc4 = 1'b1;  /* BTCLR,saddr.3,$addr8 */
                {8'h31,8'h40} : dec_pc_inc4 = 1'b1;  /* BTCLR,saddr.4,$addr8 */
                {8'h31,8'h50} : dec_pc_inc4 = 1'b1;  /* BTCLR,saddr.5,$addr8 */
                {8'h31,8'h60} : dec_pc_inc4 = 1'b1;  /* BTCLR,saddr.6,$addr8 */
                {8'h31,8'h70} : dec_pc_inc4 = 1'b1;  /* BTCLR,saddr.7,$addr8 */
                {8'h31,8'h80} : dec_pc_inc4 = 1'b1;  /* BTCLR,sfr.0,$addr8 */
                {8'h31,8'h90} : dec_pc_inc4 = 1'b1;  /* BTCLR,sfr.1,$addr8 */
                {8'h31,8'ha0} : dec_pc_inc4 = 1'b1;  /* BTCLR,sfr.2,$addr8 */
                {8'h31,8'hb0} : dec_pc_inc4 = 1'b1;  /* BTCLR,sfr.3,$addr8 */
                {8'h31,8'hc0} : dec_pc_inc4 = 1'b1;  /* BTCLR,sfr.4,$addr8 */
                {8'h31,8'hd0} : dec_pc_inc4 = 1'b1;  /* BTCLR,sfr.5,$addr8 */
                {8'h31,8'he0} : dec_pc_inc4 = 1'b1;  /* BTCLR,sfr.6,$addr8 */
                {8'h31,8'hf0} : dec_pc_inc4 = 1'b1;  /* BTCLR,sfr.7,$addr8 */
                {8'h61,8'hc1} : dec_pc_inc4 = 1'b1;  /* SOFT4,,BREAK */
                {8'h61,8'hba} : dec_pc_inc4 = 1'b1;  /* XCH,A,!addr16 */
                default : dec_pc_inc4 = 1'b0;
            endcase
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'hcf,8'hxx,2'bxx} : dec_pc_inc4 = 1'b1;  /* MOV,!addr16,#byte */
                {8'h19,8'hxx,2'bxx} : dec_pc_inc4 = 1'b1;  /* MOV,word[B],#byte */
                {8'h38,8'hxx,2'bxx} : dec_pc_inc4 = 1'b1;  /* MOV,word[C],#byte */
                {8'h39,8'hxx,2'bxx} : dec_pc_inc4 = 1'b1;  /* MOV,word[BC],#byte */
                {8'h61,8'haa,2'bx1} : dec_pc_inc4 = 1'b1;  /* XCH,A,!addr16 */
                {8'hc9,8'hxx,2'bxx} : dec_pc_inc4 = 1'b1;  /* MOVW,saddrp,#word */
                {8'hcb,8'hxx,2'bxx} : dec_pc_inc4 = 1'b1;  /* MOVW,sfrp,#word */
                {8'h40,8'hxx,2'bxx} : dec_pc_inc4 = 1'b1;  /* CMP,!addr16,#byte */
                {8'h71,8'h00,2'bx1} : dec_pc_inc4 = 1'b1;  /* SET1,,!addr16.0 */
                {8'h71,8'h10,2'bx1} : dec_pc_inc4 = 1'b1;  /* SET1,,!addr16.1 */
                {8'h71,8'h20,2'bx1} : dec_pc_inc4 = 1'b1;  /* SET1,,!addr16.2 */
                {8'h71,8'h30,2'bx1} : dec_pc_inc4 = 1'b1;  /* SET1,,!addr16.3 */
                {8'h71,8'h40,2'bx1} : dec_pc_inc4 = 1'b1;  /* SET1,,!addr16.4 */
                {8'h71,8'h50,2'bx1} : dec_pc_inc4 = 1'b1;  /* SET1,,!addr16.5 */
                {8'h71,8'h60,2'bx1} : dec_pc_inc4 = 1'b1;  /* SET1,,!addr16.6 */
                {8'h71,8'h70,2'bx1} : dec_pc_inc4 = 1'b1;  /* SET1,,!addr16.7 */
                {8'h71,8'h08,2'bx1} : dec_pc_inc4 = 1'b1;  /* CLR1,,!addr16.0 */
                {8'h71,8'h18,2'bx1} : dec_pc_inc4 = 1'b1;  /* CLR1,,!addr16.1 */
                {8'h71,8'h28,2'bx1} : dec_pc_inc4 = 1'b1;  /* CLR1,,!addr16.2 */
                {8'h71,8'h38,2'bx1} : dec_pc_inc4 = 1'b1;  /* CLR1,,!addr16.3 */
                {8'h71,8'h48,2'bx1} : dec_pc_inc4 = 1'b1;  /* CLR1,,!addr16.4 */
                {8'h71,8'h58,2'bx1} : dec_pc_inc4 = 1'b1;  /* CLR1,,!addr16.5 */
                {8'h71,8'h68,2'bx1} : dec_pc_inc4 = 1'b1;  /* CLR1,,!addr16.6 */
                {8'h71,8'h78,2'bx1} : dec_pc_inc4 = 1'b1;  /* CLR1,,!addr16.7 */
                {8'hfc,8'hxx,2'bx0} : dec_pc_inc4 = 1'b1;  /* CALL,,!!addr20 */
                {8'h31,8'h02,2'b10} : dec_pc_inc4 = 1'b1;  /* BT,saddr.0,$addr8 */
                {8'h31,8'h12,2'b10} : dec_pc_inc4 = 1'b1;  /* BT,saddr.1,$addr8 */
                {8'h31,8'h22,2'b10} : dec_pc_inc4 = 1'b1;  /* BT,saddr.2,$addr8 */
                {8'h31,8'h32,2'b10} : dec_pc_inc4 = 1'b1;  /* BT,saddr.3,$addr8 */
                {8'h31,8'h42,2'b10} : dec_pc_inc4 = 1'b1;  /* BT,saddr.4,$addr8 */
                {8'h31,8'h52,2'b10} : dec_pc_inc4 = 1'b1;  /* BT,saddr.5,$addr8 */
                {8'h31,8'h62,2'b10} : dec_pc_inc4 = 1'b1;  /* BT,saddr.6,$addr8 */
                {8'h31,8'h72,2'b10} : dec_pc_inc4 = 1'b1;  /* BT,saddr.7,$addr8 */
                {8'h31,8'h82,2'b10} : dec_pc_inc4 = 1'b1;  /* BT,sfr.0,$addr8 */
                {8'h31,8'h92,2'b10} : dec_pc_inc4 = 1'b1;  /* BT,sfr.1,$addr8 */
                {8'h31,8'ha2,2'b10} : dec_pc_inc4 = 1'b1;  /* BT,sfr.2,$addr8 */
                {8'h31,8'hb2,2'b10} : dec_pc_inc4 = 1'b1;  /* BT,sfr.3,$addr8 */
                {8'h31,8'hc2,2'b10} : dec_pc_inc4 = 1'b1;  /* BT,sfr.4,$addr8 */
                {8'h31,8'hd2,2'b10} : dec_pc_inc4 = 1'b1;  /* BT,sfr.5,$addr8 */
                {8'h31,8'he2,2'b10} : dec_pc_inc4 = 1'b1;  /* BT,sfr.6,$addr8 */
                {8'h31,8'hf2,2'b10} : dec_pc_inc4 = 1'b1;  /* BT,sfr.7,$addr8 */
                {8'h31,8'h04,2'b10} : dec_pc_inc4 = 1'b1;  /* BF,saddr.0,$addr8 */
                {8'h31,8'h14,2'b10} : dec_pc_inc4 = 1'b1;  /* BF,saddr.1,$addr8 */
                {8'h31,8'h24,2'b10} : dec_pc_inc4 = 1'b1;  /* BF,saddr.2,$addr8 */
                {8'h31,8'h34,2'b10} : dec_pc_inc4 = 1'b1;  /* BF,saddr.3,$addr8 */
                {8'h31,8'h44,2'b10} : dec_pc_inc4 = 1'b1;  /* BF,saddr.4,$addr8 */
                {8'h31,8'h54,2'b10} : dec_pc_inc4 = 1'b1;  /* BF,saddr.5,$addr8 */
                {8'h31,8'h64,2'b10} : dec_pc_inc4 = 1'b1;  /* BF,saddr.6,$addr8 */
                {8'h31,8'h74,2'b10} : dec_pc_inc4 = 1'b1;  /* BF,saddr.7,$addr8 */
                {8'h31,8'h84,2'b10} : dec_pc_inc4 = 1'b1;  /* BF,sfr.0,$addr8 */
                {8'h31,8'h94,2'b10} : dec_pc_inc4 = 1'b1;  /* BF,sfr.1,$addr8 */
                {8'h31,8'ha4,2'b10} : dec_pc_inc4 = 1'b1;  /* BF,sfr.2,$addr8 */
                {8'h31,8'hb4,2'b10} : dec_pc_inc4 = 1'b1;  /* BF,sfr.3,$addr8 */
                {8'h31,8'hc4,2'b10} : dec_pc_inc4 = 1'b1;  /* BF,sfr.4,$addr8 */
                {8'h31,8'hd4,2'b10} : dec_pc_inc4 = 1'b1;  /* BF,sfr.5,$addr8 */
                {8'h31,8'he4,2'b10} : dec_pc_inc4 = 1'b1;  /* BF,sfr.6,$addr8 */
                {8'h31,8'hf4,2'b10} : dec_pc_inc4 = 1'b1;  /* BF,sfr.7,$addr8 */
                {8'h31,8'h00,2'b10} : dec_pc_inc4 = 1'b1;  /* BTCLR,saddr.0,$addr8 */
                {8'h31,8'h10,2'b10} : dec_pc_inc4 = 1'b1;  /* BTCLR,saddr.1,$addr8 */
                {8'h31,8'h20,2'b10} : dec_pc_inc4 = 1'b1;  /* BTCLR,saddr.2,$addr8 */
                {8'h31,8'h30,2'b10} : dec_pc_inc4 = 1'b1;  /* BTCLR,saddr.3,$addr8 */
                {8'h31,8'h40,2'b10} : dec_pc_inc4 = 1'b1;  /* BTCLR,saddr.4,$addr8 */
                {8'h31,8'h50,2'b10} : dec_pc_inc4 = 1'b1;  /* BTCLR,saddr.5,$addr8 */
                {8'h31,8'h60,2'b10} : dec_pc_inc4 = 1'b1;  /* BTCLR,saddr.6,$addr8 */
                {8'h31,8'h70,2'b10} : dec_pc_inc4 = 1'b1;  /* BTCLR,saddr.7,$addr8 */
                {8'h31,8'h80,2'b10} : dec_pc_inc4 = 1'b1;  /* BTCLR,sfr.0,$addr8 */
                {8'h31,8'h90,2'b10} : dec_pc_inc4 = 1'b1;  /* BTCLR,sfr.1,$addr8 */
                {8'h31,8'ha0,2'b10} : dec_pc_inc4 = 1'b1;  /* BTCLR,sfr.2,$addr8 */
                {8'h31,8'hb0,2'b10} : dec_pc_inc4 = 1'b1;  /* BTCLR,sfr.3,$addr8 */
                {8'h31,8'hc0,2'b10} : dec_pc_inc4 = 1'b1;  /* BTCLR,sfr.4,$addr8 */
                {8'h31,8'hd0,2'b10} : dec_pc_inc4 = 1'b1;  /* BTCLR,sfr.5,$addr8 */
                {8'h31,8'he0,2'b10} : dec_pc_inc4 = 1'b1;  /* BTCLR,sfr.6,$addr8 */
                {8'h31,8'hf0,2'b10} : dec_pc_inc4 = 1'b1;  /* BTCLR,sfr.7,$addr8 */
                {8'h61,8'hc1,2'bx0} : dec_pc_inc4 = 1'b1;  /* SOFT4,,BREAK */
                {8'h61,8'hba,2'bx1} : dec_pc_inc4 = 1'b1;  /* XCH,A,!addr16 */
                default : dec_pc_inc4 = 1'b0;
            endcase
        end
    end
    output dec_clear_stage;
    reg    dec_clear_stage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1) begin
            dec_clear_stage = 1'b1;  /* RESET */
        end else if(ivack == 1'b1) begin
            casex ({stage_adr})  
                {2'b00} : dec_clear_stage = 1'b0;  /* Interrupt */
                {2'b01} : dec_clear_stage = 1'b0;  /* Interrupt */
                {2'b10} : dec_clear_stage = 1'b0;  /* Interrupt */
                default : dec_clear_stage = 1'b1;
            endcase
        end else if(skpack == 1'b1) begin
            dec_clear_stage = 1'b1;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'ha8,2'bx0} : dec_clear_stage = 1'b0;  /* XCH,A,saddr */
                {8'h61,8'hab,2'bx0} : dec_clear_stage = 1'b0;  /* XCH,A,sfr */
                {8'h61,8'haa,2'bx0} : dec_clear_stage = 1'b0;  /* XCH,A,!addr16 */
                {8'h61,8'hae,2'bx0} : dec_clear_stage = 1'b0;  /* XCH,A,[DE] */
                {8'h61,8'haf,2'bx0} : dec_clear_stage = 1'b0;  /* XCH,A,[DE+byte] */
                {8'h61,8'hac,2'bx0} : dec_clear_stage = 1'b0;  /* XCH,A,[HL] */
                {8'h61,8'had,2'bx0} : dec_clear_stage = 1'b0;  /* XCH,A,[HL+byte] */
                {8'h61,8'hb9,2'bx0} : dec_clear_stage = 1'b0;  /* XCH,A,[HL+B] */
                {8'h61,8'ha9,2'bx0} : dec_clear_stage = 1'b0;  /* XCH,A,[HL+C] */
                {8'h0a,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* ADD,saddr,#byte */
                {8'h1a,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* ADDC,saddr,#byte */
                {8'h2a,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* SUB,saddr,#byte */
                {8'h3a,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* SUBC,saddr,#byte */
                {8'h5a,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* AND,saddr,#byte */
                {8'h6a,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* OR,saddr,#byte */
                {8'h7a,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* XOR,saddr,#byte */
                {8'ha4,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* INC,,saddr */
                {8'ha0,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* INC,,!addr16 */
                {8'h61,8'h59,2'bx0} : dec_clear_stage = 1'b0;  /* INC,,[HL+byte] */
                {8'hb4,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* DEC,,saddr */
                {8'hb0,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* DEC,,!addr16 */
                {8'h61,8'h69,2'bx0} : dec_clear_stage = 1'b0;  /* DEC,,[HL+byte] */
                {8'ha6,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* INCW,,saddrp */
                {8'ha2,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* INCW,,!addr16 */
                {8'h61,8'h79,2'bx0} : dec_clear_stage = 1'b0;  /* INCW,,[HL+byte] */
                {8'hb6,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* DECW,,saddrp */
                {8'hb2,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* DECW,,!addr16 */
                {8'h61,8'h89,2'bx0} : dec_clear_stage = 1'b0;  /* DECW,,[HL+byte] */
                {8'h71,8'h01,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,saddr.0,CY */
                {8'h71,8'h11,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,saddr.1,CY */
                {8'h71,8'h21,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,saddr.2,CY */
                {8'h71,8'h31,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,saddr.3,CY */
                {8'h71,8'h41,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,saddr.4,CY */
                {8'h71,8'h51,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,saddr.5,CY */
                {8'h71,8'h61,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,saddr.6,CY */
                {8'h71,8'h71,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,saddr.7,CY */
                {8'h71,8'h09,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,sfr.0,CY */
                {8'h71,8'h19,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,sfr.1,CY */
                {8'h71,8'h29,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,sfr.2,CY */
                {8'h71,8'h39,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,sfr.3,CY */
                {8'h71,8'h49,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,sfr.4,CY */
                {8'h71,8'h59,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,sfr.5,CY */
                {8'h71,8'h69,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,sfr.6,CY */
                {8'h71,8'h79,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,sfr.7,CY */
                {8'h71,8'h81,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,[HL].0,CY */
                {8'h71,8'h91,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,[HL].1,CY */
                {8'h71,8'ha1,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,[HL].2,CY */
                {8'h71,8'hb1,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,[HL].3,CY */
                {8'h71,8'hc1,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,[HL].4,CY */
                {8'h71,8'hd1,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,[HL].5,CY */
                {8'h71,8'he1,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,[HL].6,CY */
                {8'h71,8'hf1,2'bx0} : dec_clear_stage = 1'b0;  /* MOV1,[HL].7,CY */
                {8'h71,8'h02,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,saddr.0 */
                {8'h71,8'h12,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,saddr.1 */
                {8'h71,8'h22,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,saddr.2 */
                {8'h71,8'h32,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,saddr.3 */
                {8'h71,8'h42,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,saddr.4 */
                {8'h71,8'h52,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,saddr.5 */
                {8'h71,8'h62,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,saddr.6 */
                {8'h71,8'h72,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,saddr.7 */
                {8'h71,8'h0a,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,sfr.0 */
                {8'h71,8'h1a,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,sfr.1 */
                {8'h71,8'h2a,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,sfr.2 */
                {8'h71,8'h3a,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,sfr.3 */
                {8'h71,8'h4a,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,sfr.4 */
                {8'h71,8'h5a,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,sfr.5 */
                {8'h71,8'h6a,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,sfr.6 */
                {8'h71,8'h7a,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,sfr.7 */
                {8'h71,8'h00,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,!addr16.0 */
                {8'h71,8'h10,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,!addr16.1 */
                {8'h71,8'h20,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,!addr16.2 */
                {8'h71,8'h30,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,!addr16.3 */
                {8'h71,8'h40,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,!addr16.4 */
                {8'h71,8'h50,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,!addr16.5 */
                {8'h71,8'h60,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,!addr16.6 */
                {8'h71,8'h70,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,!addr16.7 */
                {8'h71,8'h82,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,[HL].0 */
                {8'h71,8'h92,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,[HL].1 */
                {8'h71,8'ha2,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,[HL].2 */
                {8'h71,8'hb2,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,[HL].3 */
                {8'h71,8'hc2,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,[HL].4 */
                {8'h71,8'hd2,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,[HL].5 */
                {8'h71,8'he2,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,[HL].6 */
                {8'h71,8'hf2,2'bx0} : dec_clear_stage = 1'b0;  /* SET1,,[HL].7 */
                {8'h71,8'h03,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,saddr.0 */
                {8'h71,8'h13,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,saddr.1 */
                {8'h71,8'h23,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,saddr.2 */
                {8'h71,8'h33,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,saddr.3 */
                {8'h71,8'h43,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,saddr.4 */
                {8'h71,8'h53,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,saddr.5 */
                {8'h71,8'h63,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,saddr.6 */
                {8'h71,8'h73,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,saddr.7 */
                {8'h71,8'h0b,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,sfr.0 */
                {8'h71,8'h1b,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,sfr.1 */
                {8'h71,8'h2b,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,sfr.2 */
                {8'h71,8'h3b,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,sfr.3 */
                {8'h71,8'h4b,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,sfr.4 */
                {8'h71,8'h5b,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,sfr.5 */
                {8'h71,8'h6b,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,sfr.6 */
                {8'h71,8'h7b,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,sfr.7 */
                {8'h71,8'h08,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,!addr16.0 */
                {8'h71,8'h18,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,!addr16.1 */
                {8'h71,8'h28,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,!addr16.2 */
                {8'h71,8'h38,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,!addr16.3 */
                {8'h71,8'h48,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,!addr16.4 */
                {8'h71,8'h58,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,!addr16.5 */
                {8'h71,8'h68,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,!addr16.6 */
                {8'h71,8'h78,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,!addr16.7 */
                {8'h71,8'h83,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,[HL].0 */
                {8'h71,8'h93,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,[HL].1 */
                {8'h71,8'ha3,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,[HL].2 */
                {8'h71,8'hb3,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,[HL].3 */
                {8'h71,8'hc3,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,[HL].4 */
                {8'h71,8'hd3,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,[HL].5 */
                {8'h71,8'he3,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,[HL].6 */
                {8'h71,8'hf3,2'bx0} : dec_clear_stage = 1'b0;  /* CLR1,,[HL].7 */
                {8'h61,8'hca,2'bx0} : dec_clear_stage = 1'b0;  /* CALL,,AX */
                {8'h61,8'hda,2'bx0} : dec_clear_stage = 1'b0;  /* CALL,,BC */
                {8'h61,8'hea,2'bx0} : dec_clear_stage = 1'b0;  /* CALL,,DE */
                {8'h61,8'hfa,2'bx0} : dec_clear_stage = 1'b0;  /* CALL,,HL */
                {8'hfe,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* CALL,,$!addr16 */
                {8'hfd,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* CALL,,!addr16 */
                {8'hfc,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* CALL,,!!addr20 */
                {8'h61,8'h84,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[0080h] */
                {8'h61,8'h94,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[0082h] */
                {8'h61,8'ha4,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[0084h] */
                {8'h61,8'hb4,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[0086h] */
                {8'h61,8'hc4,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[0088h] */
                {8'h61,8'hd4,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[008Ah] */
                {8'h61,8'he4,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[008Ch] */
                {8'h61,8'hf4,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[008Eh] */
                {8'h61,8'h85,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[0090h] */
                {8'h61,8'h95,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[0092h] */
                {8'h61,8'ha5,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[0094h] */
                {8'h61,8'hb5,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[0096h] */
                {8'h61,8'hc5,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[0098h] */
                {8'h61,8'hd5,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[009Ah] */
                {8'h61,8'he5,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[009Ch] */
                {8'h61,8'hf5,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[009Eh] */
                {8'h61,8'h86,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[00A0h] */
                {8'h61,8'h96,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[00A2h] */
                {8'h61,8'ha6,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[00A4h] */
                {8'h61,8'hb6,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[00A6h] */
                {8'h61,8'hc6,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[00A8h] */
                {8'h61,8'hd6,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[00AAh] */
                {8'h61,8'he6,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[00ACh] */
                {8'h61,8'hf6,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[00AEh] */
                {8'h61,8'h87,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[00B0h] */
                {8'h61,8'h97,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[00B2h] */
                {8'h61,8'ha7,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[00B4h] */
                {8'h61,8'hb7,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[00B6h] */
                {8'h61,8'hc7,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[00B8h] */
                {8'h61,8'hd7,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[00BAh] */
                {8'h61,8'he7,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[00BCh] */
                {8'h61,8'hf7,2'bx0} : dec_clear_stage = 1'b0;  /* CALLT,,[00BEh] */
                {8'h61,8'hcc,2'bx0} : dec_clear_stage = 1'b0;  /* BRK,, */
                {8'hd7,8'hxx,2'b00} : dec_clear_stage = 1'b0;  /* RET,, */
                {8'hd7,8'hxx,2'b01} : dec_clear_stage = 1'b0;  /* RET,, */
                {8'hd7,8'hxx,2'b10} : dec_clear_stage = 1'b0;  /* RET,, */
                {8'h61,8'hec,2'b00} : dec_clear_stage = 1'b0;  /* RETB,, */
                {8'h61,8'hec,2'b01} : dec_clear_stage = 1'b0;  /* RETB,, */
                {8'h61,8'hec,2'b10} : dec_clear_stage = 1'b0;  /* RETB,, */
                {8'h61,8'hfc,2'b00} : dec_clear_stage = 1'b0;  /* RETI,, */
                {8'h61,8'hfc,2'b01} : dec_clear_stage = 1'b0;  /* RETI,, */
                {8'h61,8'hfc,2'b10} : dec_clear_stage = 1'b0;  /* RETI,, */
                {8'hec,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* BR,,!!addr20 */
                {8'hed,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* BR,,!addr16 */
                {8'hee,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* BR,,$!addr16 */
                {8'hef,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* BR,,$addr8 */
                {8'h61,8'hcb,2'bx0} : dec_clear_stage = 1'b0;  /* BR,,AX */
                {8'hdc,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* BC,,$addr8 */
                {8'hde,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* BNC,,$addr8 */
                {8'hdd,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* BZ,,$addr8 */
                {8'hdf,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* BNZ,,$addr8 */
                {8'h61,8'hc3,2'bx0} : dec_clear_stage = 1'b0;  /* BH,,$addr8 */
                {8'h61,8'hd3,2'bx0} : dec_clear_stage = 1'b0;  /* BNH,,$addr8 */
                {8'h31,8'h02,2'b00} : dec_clear_stage = 1'b0;  /* BT,saddr.0,$addr8 */
                {8'h31,8'h02,2'b01} : dec_clear_stage = 1'b0;  /* BT,saddr.0,$addr8 */
                {8'h31,8'h12,2'b00} : dec_clear_stage = 1'b0;  /* BT,saddr.1,$addr8 */
                {8'h31,8'h12,2'b01} : dec_clear_stage = 1'b0;  /* BT,saddr.1,$addr8 */
                {8'h31,8'h22,2'b00} : dec_clear_stage = 1'b0;  /* BT,saddr.2,$addr8 */
                {8'h31,8'h22,2'b01} : dec_clear_stage = 1'b0;  /* BT,saddr.2,$addr8 */
                {8'h31,8'h32,2'b00} : dec_clear_stage = 1'b0;  /* BT,saddr.3,$addr8 */
                {8'h31,8'h32,2'b01} : dec_clear_stage = 1'b0;  /* BT,saddr.3,$addr8 */
                {8'h31,8'h42,2'b00} : dec_clear_stage = 1'b0;  /* BT,saddr.4,$addr8 */
                {8'h31,8'h42,2'b01} : dec_clear_stage = 1'b0;  /* BT,saddr.4,$addr8 */
                {8'h31,8'h52,2'b00} : dec_clear_stage = 1'b0;  /* BT,saddr.5,$addr8 */
                {8'h31,8'h52,2'b01} : dec_clear_stage = 1'b0;  /* BT,saddr.5,$addr8 */
                {8'h31,8'h62,2'b00} : dec_clear_stage = 1'b0;  /* BT,saddr.6,$addr8 */
                {8'h31,8'h62,2'b01} : dec_clear_stage = 1'b0;  /* BT,saddr.6,$addr8 */
                {8'h31,8'h72,2'b00} : dec_clear_stage = 1'b0;  /* BT,saddr.7,$addr8 */
                {8'h31,8'h72,2'b01} : dec_clear_stage = 1'b0;  /* BT,saddr.7,$addr8 */
                {8'h31,8'h82,2'b00} : dec_clear_stage = 1'b0;  /* BT,sfr.0,$addr8 */
                {8'h31,8'h82,2'b01} : dec_clear_stage = 1'b0;  /* BT,sfr.0,$addr8 */
                {8'h31,8'h92,2'b00} : dec_clear_stage = 1'b0;  /* BT,sfr.1,$addr8 */
                {8'h31,8'h92,2'b01} : dec_clear_stage = 1'b0;  /* BT,sfr.1,$addr8 */
                {8'h31,8'ha2,2'b00} : dec_clear_stage = 1'b0;  /* BT,sfr.2,$addr8 */
                {8'h31,8'ha2,2'b01} : dec_clear_stage = 1'b0;  /* BT,sfr.2,$addr8 */
                {8'h31,8'hb2,2'b00} : dec_clear_stage = 1'b0;  /* BT,sfr.3,$addr8 */
                {8'h31,8'hb2,2'b01} : dec_clear_stage = 1'b0;  /* BT,sfr.3,$addr8 */
                {8'h31,8'hc2,2'b00} : dec_clear_stage = 1'b0;  /* BT,sfr.4,$addr8 */
                {8'h31,8'hc2,2'b01} : dec_clear_stage = 1'b0;  /* BT,sfr.4,$addr8 */
                {8'h31,8'hd2,2'b00} : dec_clear_stage = 1'b0;  /* BT,sfr.5,$addr8 */
                {8'h31,8'hd2,2'b01} : dec_clear_stage = 1'b0;  /* BT,sfr.5,$addr8 */
                {8'h31,8'he2,2'b00} : dec_clear_stage = 1'b0;  /* BT,sfr.6,$addr8 */
                {8'h31,8'he2,2'b01} : dec_clear_stage = 1'b0;  /* BT,sfr.6,$addr8 */
                {8'h31,8'hf2,2'b00} : dec_clear_stage = 1'b0;  /* BT,sfr.7,$addr8 */
                {8'h31,8'hf2,2'b01} : dec_clear_stage = 1'b0;  /* BT,sfr.7,$addr8 */
                {8'h31,8'h03,2'b00} : dec_clear_stage = 1'b0;  /* BT,A.0,$addr8 */
                {8'h31,8'h03,2'b01} : dec_clear_stage = 1'b0;  /* BT,A.0,$addr8 */
                {8'h31,8'h13,2'b00} : dec_clear_stage = 1'b0;  /* BT,A.1,$addr8 */
                {8'h31,8'h13,2'b01} : dec_clear_stage = 1'b0;  /* BT,A.1,$addr8 */
                {8'h31,8'h23,2'b00} : dec_clear_stage = 1'b0;  /* BT,A.2,$addr8 */
                {8'h31,8'h23,2'b01} : dec_clear_stage = 1'b0;  /* BT,A.2,$addr8 */
                {8'h31,8'h33,2'b00} : dec_clear_stage = 1'b0;  /* BT,A.3,$addr8 */
                {8'h31,8'h33,2'b01} : dec_clear_stage = 1'b0;  /* BT,A.3,$addr8 */
                {8'h31,8'h43,2'b00} : dec_clear_stage = 1'b0;  /* BT,A.4,$addr8 */
                {8'h31,8'h43,2'b01} : dec_clear_stage = 1'b0;  /* BT,A.4,$addr8 */
                {8'h31,8'h53,2'b00} : dec_clear_stage = 1'b0;  /* BT,A.5,$addr8 */
                {8'h31,8'h53,2'b01} : dec_clear_stage = 1'b0;  /* BT,A.5,$addr8 */
                {8'h31,8'h63,2'b00} : dec_clear_stage = 1'b0;  /* BT,A.6,$addr8 */
                {8'h31,8'h63,2'b01} : dec_clear_stage = 1'b0;  /* BT,A.6,$addr8 */
                {8'h31,8'h73,2'b00} : dec_clear_stage = 1'b0;  /* BT,A.7,$addr8 */
                {8'h31,8'h73,2'b01} : dec_clear_stage = 1'b0;  /* BT,A.7,$addr8 */
                {8'h31,8'h83,2'b00} : dec_clear_stage = 1'b0;  /* BT,[HL].0,$addr8 */
                {8'h31,8'h83,2'b01} : dec_clear_stage = 1'b0;  /* BT,[HL].0,$addr8 */
                {8'h31,8'h93,2'b00} : dec_clear_stage = 1'b0;  /* BT,[HL].1,$addr8 */
                {8'h31,8'h93,2'b01} : dec_clear_stage = 1'b0;  /* BT,[HL].1,$addr8 */
                {8'h31,8'ha3,2'b00} : dec_clear_stage = 1'b0;  /* BT,[HL].2,$addr8 */
                {8'h31,8'ha3,2'b01} : dec_clear_stage = 1'b0;  /* BT,[HL].2,$addr8 */
                {8'h31,8'hb3,2'b00} : dec_clear_stage = 1'b0;  /* BT,[HL].3,$addr8 */
                {8'h31,8'hb3,2'b01} : dec_clear_stage = 1'b0;  /* BT,[HL].3,$addr8 */
                {8'h31,8'hc3,2'b00} : dec_clear_stage = 1'b0;  /* BT,[HL].4,$addr8 */
                {8'h31,8'hc3,2'b01} : dec_clear_stage = 1'b0;  /* BT,[HL].4,$addr8 */
                {8'h31,8'hd3,2'b00} : dec_clear_stage = 1'b0;  /* BT,[HL].5,$addr8 */
                {8'h31,8'hd3,2'b01} : dec_clear_stage = 1'b0;  /* BT,[HL].5,$addr8 */
                {8'h31,8'he3,2'b00} : dec_clear_stage = 1'b0;  /* BT,[HL].6,$addr8 */
                {8'h31,8'he3,2'b01} : dec_clear_stage = 1'b0;  /* BT,[HL].6,$addr8 */
                {8'h31,8'hf3,2'b00} : dec_clear_stage = 1'b0;  /* BT,[HL].7,$addr8 */
                {8'h31,8'hf3,2'b01} : dec_clear_stage = 1'b0;  /* BT,[HL].7,$addr8 */
                {8'h31,8'h04,2'b00} : dec_clear_stage = 1'b0;  /* BF,saddr.0,$addr8 */
                {8'h31,8'h04,2'b01} : dec_clear_stage = 1'b0;  /* BF,saddr.0,$addr8 */
                {8'h31,8'h14,2'b00} : dec_clear_stage = 1'b0;  /* BF,saddr.1,$addr8 */
                {8'h31,8'h14,2'b01} : dec_clear_stage = 1'b0;  /* BF,saddr.1,$addr8 */
                {8'h31,8'h24,2'b00} : dec_clear_stage = 1'b0;  /* BF,saddr.2,$addr8 */
                {8'h31,8'h24,2'b01} : dec_clear_stage = 1'b0;  /* BF,saddr.2,$addr8 */
                {8'h31,8'h34,2'b00} : dec_clear_stage = 1'b0;  /* BF,saddr.3,$addr8 */
                {8'h31,8'h34,2'b01} : dec_clear_stage = 1'b0;  /* BF,saddr.3,$addr8 */
                {8'h31,8'h44,2'b00} : dec_clear_stage = 1'b0;  /* BF,saddr.4,$addr8 */
                {8'h31,8'h44,2'b01} : dec_clear_stage = 1'b0;  /* BF,saddr.4,$addr8 */
                {8'h31,8'h54,2'b00} : dec_clear_stage = 1'b0;  /* BF,saddr.5,$addr8 */
                {8'h31,8'h54,2'b01} : dec_clear_stage = 1'b0;  /* BF,saddr.5,$addr8 */
                {8'h31,8'h64,2'b00} : dec_clear_stage = 1'b0;  /* BF,saddr.6,$addr8 */
                {8'h31,8'h64,2'b01} : dec_clear_stage = 1'b0;  /* BF,saddr.6,$addr8 */
                {8'h31,8'h74,2'b00} : dec_clear_stage = 1'b0;  /* BF,saddr.7,$addr8 */
                {8'h31,8'h74,2'b01} : dec_clear_stage = 1'b0;  /* BF,saddr.7,$addr8 */
                {8'h31,8'h84,2'b00} : dec_clear_stage = 1'b0;  /* BF,sfr.0,$addr8 */
                {8'h31,8'h84,2'b01} : dec_clear_stage = 1'b0;  /* BF,sfr.0,$addr8 */
                {8'h31,8'h94,2'b00} : dec_clear_stage = 1'b0;  /* BF,sfr.1,$addr8 */
                {8'h31,8'h94,2'b01} : dec_clear_stage = 1'b0;  /* BF,sfr.1,$addr8 */
                {8'h31,8'ha4,2'b00} : dec_clear_stage = 1'b0;  /* BF,sfr.2,$addr8 */
                {8'h31,8'ha4,2'b01} : dec_clear_stage = 1'b0;  /* BF,sfr.2,$addr8 */
                {8'h31,8'hb4,2'b00} : dec_clear_stage = 1'b0;  /* BF,sfr.3,$addr8 */
                {8'h31,8'hb4,2'b01} : dec_clear_stage = 1'b0;  /* BF,sfr.3,$addr8 */
                {8'h31,8'hc4,2'b00} : dec_clear_stage = 1'b0;  /* BF,sfr.4,$addr8 */
                {8'h31,8'hc4,2'b01} : dec_clear_stage = 1'b0;  /* BF,sfr.4,$addr8 */
                {8'h31,8'hd4,2'b00} : dec_clear_stage = 1'b0;  /* BF,sfr.5,$addr8 */
                {8'h31,8'hd4,2'b01} : dec_clear_stage = 1'b0;  /* BF,sfr.5,$addr8 */
                {8'h31,8'he4,2'b00} : dec_clear_stage = 1'b0;  /* BF,sfr.6,$addr8 */
                {8'h31,8'he4,2'b01} : dec_clear_stage = 1'b0;  /* BF,sfr.6,$addr8 */
                {8'h31,8'hf4,2'b00} : dec_clear_stage = 1'b0;  /* BF,sfr.7,$addr8 */
                {8'h31,8'hf4,2'b01} : dec_clear_stage = 1'b0;  /* BF,sfr.7,$addr8 */
                {8'h31,8'h05,2'b00} : dec_clear_stage = 1'b0;  /* BF,A.0,$addr8 */
                {8'h31,8'h05,2'b01} : dec_clear_stage = 1'b0;  /* BF,A.0,$addr8 */
                {8'h31,8'h15,2'b00} : dec_clear_stage = 1'b0;  /* BF,A.1,$addr8 */
                {8'h31,8'h15,2'b01} : dec_clear_stage = 1'b0;  /* BF,A.1,$addr8 */
                {8'h31,8'h25,2'b00} : dec_clear_stage = 1'b0;  /* BF,A.2,$addr8 */
                {8'h31,8'h25,2'b01} : dec_clear_stage = 1'b0;  /* BF,A.2,$addr8 */
                {8'h31,8'h35,2'b00} : dec_clear_stage = 1'b0;  /* BF,A.3,$addr8 */
                {8'h31,8'h35,2'b01} : dec_clear_stage = 1'b0;  /* BF,A.3,$addr8 */
                {8'h31,8'h45,2'b00} : dec_clear_stage = 1'b0;  /* BF,A.4,$addr8 */
                {8'h31,8'h45,2'b01} : dec_clear_stage = 1'b0;  /* BF,A.4,$addr8 */
                {8'h31,8'h55,2'b00} : dec_clear_stage = 1'b0;  /* BF,A.5,$addr8 */
                {8'h31,8'h55,2'b01} : dec_clear_stage = 1'b0;  /* BF,A.5,$addr8 */
                {8'h31,8'h65,2'b00} : dec_clear_stage = 1'b0;  /* BF,A.6,$addr8 */
                {8'h31,8'h65,2'b01} : dec_clear_stage = 1'b0;  /* BF,A.6,$addr8 */
                {8'h31,8'h75,2'b00} : dec_clear_stage = 1'b0;  /* BF,A.7,$addr8 */
                {8'h31,8'h75,2'b01} : dec_clear_stage = 1'b0;  /* BF,A.7,$addr8 */
                {8'h31,8'h85,2'b00} : dec_clear_stage = 1'b0;  /* BF,[HL].0,$addr8 */
                {8'h31,8'h85,2'b01} : dec_clear_stage = 1'b0;  /* BF,[HL].0,$addr8 */
                {8'h31,8'h95,2'b00} : dec_clear_stage = 1'b0;  /* BF,[HL].1,$addr8 */
                {8'h31,8'h95,2'b01} : dec_clear_stage = 1'b0;  /* BF,[HL].1,$addr8 */
                {8'h31,8'ha5,2'b00} : dec_clear_stage = 1'b0;  /* BF,[HL].2,$addr8 */
                {8'h31,8'ha5,2'b01} : dec_clear_stage = 1'b0;  /* BF,[HL].2,$addr8 */
                {8'h31,8'hb5,2'b00} : dec_clear_stage = 1'b0;  /* BF,[HL].3,$addr8 */
                {8'h31,8'hb5,2'b01} : dec_clear_stage = 1'b0;  /* BF,[HL].3,$addr8 */
                {8'h31,8'hc5,2'b00} : dec_clear_stage = 1'b0;  /* BF,[HL].4,$addr8 */
                {8'h31,8'hc5,2'b01} : dec_clear_stage = 1'b0;  /* BF,[HL].4,$addr8 */
                {8'h31,8'hd5,2'b00} : dec_clear_stage = 1'b0;  /* BF,[HL].5,$addr8 */
                {8'h31,8'hd5,2'b01} : dec_clear_stage = 1'b0;  /* BF,[HL].5,$addr8 */
                {8'h31,8'he5,2'b00} : dec_clear_stage = 1'b0;  /* BF,[HL].6,$addr8 */
                {8'h31,8'he5,2'b01} : dec_clear_stage = 1'b0;  /* BF,[HL].6,$addr8 */
                {8'h31,8'hf5,2'b00} : dec_clear_stage = 1'b0;  /* BF,[HL].7,$addr8 */
                {8'h31,8'hf5,2'b01} : dec_clear_stage = 1'b0;  /* BF,[HL].7,$addr8 */
                {8'h31,8'h00,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,saddr.0,$addr8 */
                {8'h31,8'h00,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,saddr.0,$addr8 */
                {8'h31,8'h10,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,saddr.1,$addr8 */
                {8'h31,8'h10,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,saddr.1,$addr8 */
                {8'h31,8'h20,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,saddr.2,$addr8 */
                {8'h31,8'h20,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,saddr.2,$addr8 */
                {8'h31,8'h30,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,saddr.3,$addr8 */
                {8'h31,8'h30,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,saddr.3,$addr8 */
                {8'h31,8'h40,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,saddr.4,$addr8 */
                {8'h31,8'h40,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,saddr.4,$addr8 */
                {8'h31,8'h50,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,saddr.5,$addr8 */
                {8'h31,8'h50,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,saddr.5,$addr8 */
                {8'h31,8'h60,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,saddr.6,$addr8 */
                {8'h31,8'h60,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,saddr.6,$addr8 */
                {8'h31,8'h70,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,saddr.7,$addr8 */
                {8'h31,8'h70,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,saddr.7,$addr8 */
                {8'h31,8'h80,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,sfr.0,$addr8 */
                {8'h31,8'h80,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,sfr.0,$addr8 */
                {8'h31,8'h90,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,sfr.1,$addr8 */
                {8'h31,8'h90,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,sfr.1,$addr8 */
                {8'h31,8'ha0,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,sfr.2,$addr8 */
                {8'h31,8'ha0,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,sfr.2,$addr8 */
                {8'h31,8'hb0,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,sfr.3,$addr8 */
                {8'h31,8'hb0,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,sfr.3,$addr8 */
                {8'h31,8'hc0,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,sfr.4,$addr8 */
                {8'h31,8'hc0,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,sfr.4,$addr8 */
                {8'h31,8'hd0,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,sfr.5,$addr8 */
                {8'h31,8'hd0,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,sfr.5,$addr8 */
                {8'h31,8'he0,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,sfr.6,$addr8 */
                {8'h31,8'he0,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,sfr.6,$addr8 */
                {8'h31,8'hf0,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,sfr.7,$addr8 */
                {8'h31,8'hf0,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,sfr.7,$addr8 */
                {8'h31,8'h01,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,A.0,$addr8 */
                {8'h31,8'h01,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,A.0,$addr8 */
                {8'h31,8'h11,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,A.1,$addr8 */
                {8'h31,8'h11,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,A.1,$addr8 */
                {8'h31,8'h21,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,A.2,$addr8 */
                {8'h31,8'h21,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,A.2,$addr8 */
                {8'h31,8'h31,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,A.3,$addr8 */
                {8'h31,8'h31,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,A.3,$addr8 */
                {8'h31,8'h41,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,A.4,$addr8 */
                {8'h31,8'h41,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,A.4,$addr8 */
                {8'h31,8'h51,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,A.5,$addr8 */
                {8'h31,8'h51,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,A.5,$addr8 */
                {8'h31,8'h61,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,A.6,$addr8 */
                {8'h31,8'h61,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,A.6,$addr8 */
                {8'h31,8'h71,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,A.7,$addr8 */
                {8'h31,8'h71,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,A.7,$addr8 */
                {8'h31,8'h81,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,[HL].0,$addr8 */
                {8'h31,8'h81,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,[HL].0,$addr8 */
                {8'h31,8'h91,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,[HL].1,$addr8 */
                {8'h31,8'h91,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,[HL].1,$addr8 */
                {8'h31,8'ha1,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,[HL].2,$addr8 */
                {8'h31,8'ha1,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,[HL].2,$addr8 */
                {8'h31,8'hb1,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,[HL].3,$addr8 */
                {8'h31,8'hb1,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,[HL].3,$addr8 */
                {8'h31,8'hc1,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,[HL].4,$addr8 */
                {8'h31,8'hc1,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,[HL].4,$addr8 */
                {8'h31,8'hd1,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,[HL].5,$addr8 */
                {8'h31,8'hd1,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,[HL].5,$addr8 */
                {8'h31,8'he1,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,[HL].6,$addr8 */
                {8'h31,8'he1,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,[HL].6,$addr8 */
                {8'h31,8'hf1,2'b00} : dec_clear_stage = 1'b0;  /* BTCLR,[HL].7,$addr8 */
                {8'h31,8'hf1,2'b01} : dec_clear_stage = 1'b0;  /* BTCLR,[HL].7,$addr8 */
                {8'h61,8'hed,2'b00} : dec_clear_stage = 1'b0;  /* HALT,, */
                {8'h61,8'hed,2'b01} : dec_clear_stage = 1'b0;  /* HALT,, */
                {8'h61,8'hfd,2'b00} : dec_clear_stage = 1'b0;  /* STOP,, */
                {8'h61,8'hfd,2'b01} : dec_clear_stage = 1'b0;  /* STOP,, */
                {8'hff,8'hxx,2'bx0} : dec_clear_stage = 1'b0;  /* SOFT,,BREAK */
                {8'h61,8'ha1,2'bx0} : dec_clear_stage = 1'b0;  /* SOFT2,,BREAK */
                {8'h61,8'hb1,2'bx0} : dec_clear_stage = 1'b0;  /* SOFT3,,BREAK */
                {8'h61,8'hc1,2'bx0} : dec_clear_stage = 1'b0;  /* SOFT4,,BREAK */
                {8'h61,8'hbb,2'bx0} : dec_clear_stage = 1'b0;  /* XCH,A,sfr */
                {8'h61,8'hba,2'bx0} : dec_clear_stage = 1'b0;  /* XCH,A,!addr16 */
                {8'h61,8'hbe,2'bx0} : dec_clear_stage = 1'b0;  /* XCH,A,[DE] */
                {8'h61,8'hbf,2'bx0} : dec_clear_stage = 1'b0;  /* XCH,A,[DE+byte] */
                {8'h61,8'hbc,2'bx0} : dec_clear_stage = 1'b0;  /* XCH,A,[HL] */
                {8'h61,8'hbd,2'bx0} : dec_clear_stage = 1'b0;  /* XCH,A,[HL+byte] */
                default : dec_clear_stage = 1'b1;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_pc_set_enable;
    reg    dec_pc_set_enable;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1) begin
            dec_pc_set_enable = 1'b1;  /* RESET */
        end else if(ivack == 1'b1) begin
            casex ({stage_adr})  
                {2'b01} : dec_pc_set_enable = 1'b1;  /* Interrupt */
                {2'b10} : dec_pc_set_enable = 1'b1;  /* Interrupt */
                default : dec_pc_set_enable = 1'b0;
            endcase
//        end else if(skpack == 1'b1 || decout_mask == 1'b1) begin
        end else if(skpack == 1'b1) begin
            dec_pc_set_enable = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hca,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALL,,AX */
                {8'h61,8'hda,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALL,,BC */
                {8'h61,8'hea,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALL,,DE */
                {8'h61,8'hfa,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALL,,HL */
                {8'hfe,8'hxx,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALL,,$!addr16 */
                {8'hfd,8'hxx,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALL,,!addr16 */
                {8'hfc,8'hxx,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALL,,!!addr20 */
                {8'h61,8'h84,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[0080h] */
                {8'h61,8'h84,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[0080h] */
                {8'h61,8'h94,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[0082h] */
                {8'h61,8'h94,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[0082h] */
                {8'h61,8'ha4,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[0084h] */
                {8'h61,8'ha4,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[0084h] */
                {8'h61,8'hb4,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[0086h] */
                {8'h61,8'hb4,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[0086h] */
                {8'h61,8'hc4,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[0088h] */
                {8'h61,8'hc4,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[0088h] */
                {8'h61,8'hd4,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[008Ah] */
                {8'h61,8'hd4,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[008Ah] */
                {8'h61,8'he4,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[008Ch] */
                {8'h61,8'he4,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[008Ch] */
                {8'h61,8'hf4,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[008Eh] */
                {8'h61,8'hf4,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[008Eh] */
                {8'h61,8'h85,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[0090h] */
                {8'h61,8'h85,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[0090h] */
                {8'h61,8'h95,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[0092h] */
                {8'h61,8'h95,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[0092h] */
                {8'h61,8'ha5,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[0094h] */
                {8'h61,8'ha5,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[0094h] */
                {8'h61,8'hb5,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[0096h] */
                {8'h61,8'hb5,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[0096h] */
                {8'h61,8'hc5,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[0098h] */
                {8'h61,8'hc5,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[0098h] */
                {8'h61,8'hd5,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[009Ah] */
                {8'h61,8'hd5,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[009Ah] */
                {8'h61,8'he5,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[009Ch] */
                {8'h61,8'he5,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[009Ch] */
                {8'h61,8'hf5,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[009Eh] */
                {8'h61,8'hf5,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[009Eh] */
                {8'h61,8'h86,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00A0h] */
                {8'h61,8'h86,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00A0h] */
                {8'h61,8'h96,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00A2h] */
                {8'h61,8'h96,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00A2h] */
                {8'h61,8'ha6,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00A4h] */
                {8'h61,8'ha6,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00A4h] */
                {8'h61,8'hb6,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00A6h] */
                {8'h61,8'hb6,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00A6h] */
                {8'h61,8'hc6,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00A8h] */
                {8'h61,8'hc6,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00A8h] */
                {8'h61,8'hd6,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00AAh] */
                {8'h61,8'hd6,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00AAh] */
                {8'h61,8'he6,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00ACh] */
                {8'h61,8'he6,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00ACh] */
                {8'h61,8'hf6,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00AEh] */
                {8'h61,8'hf6,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00AEh] */
                {8'h61,8'h87,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00B0h] */
                {8'h61,8'h87,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00B0h] */
                {8'h61,8'h97,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00B2h] */
                {8'h61,8'h97,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00B2h] */
                {8'h61,8'ha7,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00B4h] */
                {8'h61,8'ha7,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00B4h] */
                {8'h61,8'hb7,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00B6h] */
                {8'h61,8'hb7,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00B6h] */
                {8'h61,8'hc7,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00B8h] */
                {8'h61,8'hc7,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00B8h] */
                {8'h61,8'hd7,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00BAh] */
                {8'h61,8'hd7,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00BAh] */
                {8'h61,8'he7,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00BCh] */
                {8'h61,8'he7,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00BCh] */
                {8'h61,8'hf7,2'bx0} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00BEh] */
                {8'h61,8'hf7,2'bx1} : dec_pc_set_enable = 1'b1;  /* CALLT,,[00BEh] */
                {8'h61,8'hcc,2'bx0} : dec_pc_set_enable = 1'b1;  /* BRK,, */
                {8'h61,8'hcc,2'bx1} : dec_pc_set_enable = 1'b1;  /* BRK,, */
                {8'hd7,8'hxx,2'b11} : dec_pc_set_enable = 1'b1;  /* RET,, */
                {8'h61,8'hec,2'b11} : dec_pc_set_enable = 1'b1;  /* RETB,, */
                {8'h61,8'hfc,2'b11} : dec_pc_set_enable = 1'b1;  /* RETI,, */
                {8'hec,8'hxx,2'bx0} : dec_pc_set_enable = 1'b1;  /* BR,,!!addr20 */
                {8'hed,8'hxx,2'bx0} : dec_pc_set_enable = 1'b1;  /* BR,,!addr16 */
                {8'hee,8'hxx,2'bx0} : dec_pc_set_enable = 1'b1;  /* BR,,$!addr16 */
                {8'hef,8'hxx,2'bx0} : dec_pc_set_enable = 1'b1;  /* BR,,$addr8 */
                {8'h61,8'hcb,2'bx0} : dec_pc_set_enable = 1'b1;  /* BR,,AX */
                {8'hdc,8'hxx,2'bx1} : dec_pc_set_enable = 1'b1;  /* BC,,$addr8 */
                {8'hde,8'hxx,2'bx1} : dec_pc_set_enable = 1'b1;  /* BNC,,$addr8 */
                {8'hdd,8'hxx,2'bx1} : dec_pc_set_enable = 1'b1;  /* BZ,,$addr8 */
                {8'hdf,8'hxx,2'bx1} : dec_pc_set_enable = 1'b1;  /* BNZ,,$addr8 */
                {8'h61,8'hc3,2'bx1} : dec_pc_set_enable = 1'b1;  /* BH,,$addr8 */
                {8'h61,8'hd3,2'bx1} : dec_pc_set_enable = 1'b1;  /* BNH,,$addr8 */
                {8'h31,8'h02,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,saddr.0,$addr8 */
                {8'h31,8'h12,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,saddr.1,$addr8 */
                {8'h31,8'h22,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,saddr.2,$addr8 */
                {8'h31,8'h32,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,saddr.3,$addr8 */
                {8'h31,8'h42,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,saddr.4,$addr8 */
                {8'h31,8'h52,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,saddr.5,$addr8 */
                {8'h31,8'h62,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,saddr.6,$addr8 */
                {8'h31,8'h72,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,saddr.7,$addr8 */
                {8'h31,8'h82,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,sfr.0,$addr8 */
                {8'h31,8'h92,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,sfr.1,$addr8 */
                {8'h31,8'ha2,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,sfr.2,$addr8 */
                {8'h31,8'hb2,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,sfr.3,$addr8 */
                {8'h31,8'hc2,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,sfr.4,$addr8 */
                {8'h31,8'hd2,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,sfr.5,$addr8 */
                {8'h31,8'he2,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,sfr.6,$addr8 */
                {8'h31,8'hf2,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,sfr.7,$addr8 */
                {8'h31,8'h03,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,A.0,$addr8 */
                {8'h31,8'h13,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,A.1,$addr8 */
                {8'h31,8'h23,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,A.2,$addr8 */
                {8'h31,8'h33,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,A.3,$addr8 */
                {8'h31,8'h43,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,A.4,$addr8 */
                {8'h31,8'h53,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,A.5,$addr8 */
                {8'h31,8'h63,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,A.6,$addr8 */
                {8'h31,8'h73,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,A.7,$addr8 */
                {8'h31,8'h83,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,[HL].0,$addr8 */
                {8'h31,8'h93,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,[HL].1,$addr8 */
                {8'h31,8'ha3,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,[HL].2,$addr8 */
                {8'h31,8'hb3,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,[HL].3,$addr8 */
                {8'h31,8'hc3,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,[HL].4,$addr8 */
                {8'h31,8'hd3,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,[HL].5,$addr8 */
                {8'h31,8'he3,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,[HL].6,$addr8 */
                {8'h31,8'hf3,2'b10} : dec_pc_set_enable = 1'b1;  /* BT,[HL].7,$addr8 */
                {8'h31,8'h04,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,saddr.0,$addr8 */
                {8'h31,8'h14,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,saddr.1,$addr8 */
                {8'h31,8'h24,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,saddr.2,$addr8 */
                {8'h31,8'h34,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,saddr.3,$addr8 */
                {8'h31,8'h44,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,saddr.4,$addr8 */
                {8'h31,8'h54,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,saddr.5,$addr8 */
                {8'h31,8'h64,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,saddr.6,$addr8 */
                {8'h31,8'h74,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,saddr.7,$addr8 */
                {8'h31,8'h84,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,sfr.0,$addr8 */
                {8'h31,8'h94,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,sfr.1,$addr8 */
                {8'h31,8'ha4,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,sfr.2,$addr8 */
                {8'h31,8'hb4,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,sfr.3,$addr8 */
                {8'h31,8'hc4,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,sfr.4,$addr8 */
                {8'h31,8'hd4,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,sfr.5,$addr8 */
                {8'h31,8'he4,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,sfr.6,$addr8 */
                {8'h31,8'hf4,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,sfr.7,$addr8 */
                {8'h31,8'h05,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,A.0,$addr8 */
                {8'h31,8'h15,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,A.1,$addr8 */
                {8'h31,8'h25,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,A.2,$addr8 */
                {8'h31,8'h35,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,A.3,$addr8 */
                {8'h31,8'h45,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,A.4,$addr8 */
                {8'h31,8'h55,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,A.5,$addr8 */
                {8'h31,8'h65,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,A.6,$addr8 */
                {8'h31,8'h75,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,A.7,$addr8 */
                {8'h31,8'h85,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,[HL].0,$addr8 */
                {8'h31,8'h95,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,[HL].1,$addr8 */
                {8'h31,8'ha5,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,[HL].2,$addr8 */
                {8'h31,8'hb5,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,[HL].3,$addr8 */
                {8'h31,8'hc5,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,[HL].4,$addr8 */
                {8'h31,8'hd5,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,[HL].5,$addr8 */
                {8'h31,8'he5,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,[HL].6,$addr8 */
                {8'h31,8'hf5,2'b10} : dec_pc_set_enable = 1'b1;  /* BF,[HL].7,$addr8 */
                {8'h31,8'h00,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,saddr.0,$addr8 */
                {8'h31,8'h10,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,saddr.1,$addr8 */
                {8'h31,8'h20,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,saddr.2,$addr8 */
                {8'h31,8'h30,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,saddr.3,$addr8 */
                {8'h31,8'h40,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,saddr.4,$addr8 */
                {8'h31,8'h50,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,saddr.5,$addr8 */
                {8'h31,8'h60,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,saddr.6,$addr8 */
                {8'h31,8'h70,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,saddr.7,$addr8 */
                {8'h31,8'h80,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,sfr.0,$addr8 */
                {8'h31,8'h90,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,sfr.1,$addr8 */
                {8'h31,8'ha0,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,sfr.2,$addr8 */
                {8'h31,8'hb0,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,sfr.3,$addr8 */
                {8'h31,8'hc0,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,sfr.4,$addr8 */
                {8'h31,8'hd0,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,sfr.5,$addr8 */
                {8'h31,8'he0,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,sfr.6,$addr8 */
                {8'h31,8'hf0,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,sfr.7,$addr8 */
                {8'h31,8'h01,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,A.0,$addr8 */
                {8'h31,8'h11,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,A.1,$addr8 */
                {8'h31,8'h21,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,A.2,$addr8 */
                {8'h31,8'h31,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,A.3,$addr8 */
                {8'h31,8'h41,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,A.4,$addr8 */
                {8'h31,8'h51,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,A.5,$addr8 */
                {8'h31,8'h61,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,A.6,$addr8 */
                {8'h31,8'h71,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,A.7,$addr8 */
                {8'h31,8'h81,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,[HL].0,$addr8 */
                {8'h31,8'h91,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,[HL].1,$addr8 */
                {8'h31,8'ha1,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,[HL].2,$addr8 */
                {8'h31,8'hb1,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,[HL].3,$addr8 */
                {8'h31,8'hc1,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,[HL].4,$addr8 */
                {8'h31,8'hd1,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,[HL].5,$addr8 */
                {8'h31,8'he1,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,[HL].6,$addr8 */
                {8'h31,8'hf1,2'b10} : dec_pc_set_enable = 1'b1;  /* BTCLR,[HL].7,$addr8 */
                {8'hff,8'hxx,2'bx0} : dec_pc_set_enable = 1'b1;  /* SOFT,,BREAK */
                {8'hff,8'hxx,2'bx1} : dec_pc_set_enable = 1'b1;  /* SOFT,,BREAK */
                {8'h61,8'ha1,2'bx0} : dec_pc_set_enable = 1'b1;  /* SOFT2,,BREAK */
                {8'h61,8'ha1,2'bx1} : dec_pc_set_enable = 1'b1;  /* SOFT2,,BREAK */
                {8'h61,8'hb1,2'bx0} : dec_pc_set_enable = 1'b1;  /* SOFT3,,BREAK */
                {8'h61,8'hb1,2'bx1} : dec_pc_set_enable = 1'b1;  /* SOFT3,,BREAK */
                {8'h61,8'hc1,2'bx0} : dec_pc_set_enable = 1'b1;  /* SOFT4,,BREAK */
                {8'h61,8'hc1,2'bx1} : dec_pc_set_enable = 1'b1;  /* SOFT4,,BREAK */
                default : dec_pc_set_enable = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_pc_set_op01;
    reg    dec_pc_set_op01;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1) begin
            dec_pc_set_op01 = 1'b1;  /* RESET */
        end else if(ivack == 1'b1) begin
            casex ({stage_adr})  
                {2'b10} : dec_pc_set_op01 = 1'b1;  /* Interrupt */
                default : dec_pc_set_op01 = 1'b0;
            endcase
//        end else if(skpack == 1'b1 || decout_mask == 1'b1) begin
        end else if(skpack == 1'b1) begin
            dec_pc_set_op01 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'h84,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[0080h] */
                {8'h61,8'h94,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[0082h] */
                {8'h61,8'ha4,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[0084h] */
                {8'h61,8'hb4,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[0086h] */
                {8'h61,8'hc4,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[0088h] */
                {8'h61,8'hd4,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[008Ah] */
                {8'h61,8'he4,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[008Ch] */
                {8'h61,8'hf4,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[008Eh] */
                {8'h61,8'h85,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[0090h] */
                {8'h61,8'h95,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[0092h] */
                {8'h61,8'ha5,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[0094h] */
                {8'h61,8'hb5,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[0096h] */
                {8'h61,8'hc5,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[0098h] */
                {8'h61,8'hd5,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[009Ah] */
                {8'h61,8'he5,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[009Ch] */
                {8'h61,8'hf5,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[009Eh] */
                {8'h61,8'h86,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[00A0h] */
                {8'h61,8'h96,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[00A2h] */
                {8'h61,8'ha6,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[00A4h] */
                {8'h61,8'hb6,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[00A6h] */
                {8'h61,8'hc6,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[00A8h] */
                {8'h61,8'hd6,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[00AAh] */
                {8'h61,8'he6,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[00ACh] */
                {8'h61,8'hf6,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[00AEh] */
                {8'h61,8'h87,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[00B0h] */
                {8'h61,8'h97,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[00B2h] */
                {8'h61,8'ha7,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[00B4h] */
                {8'h61,8'hb7,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[00B6h] */
                {8'h61,8'hc7,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[00B8h] */
                {8'h61,8'hd7,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[00BAh] */
                {8'h61,8'he7,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[00BCh] */
                {8'h61,8'hf7,2'bx1} : dec_pc_set_op01 = 1'b1;  /* CALLT,,[00BEh] */
                {8'h61,8'hcc,2'bx1} : dec_pc_set_op01 = 1'b1;  /* BRK,, */
                {8'hff,8'hxx,2'bx1} : dec_pc_set_op01 = 1'b1;  /* SOFT,,BREAK */
                {8'h61,8'ha1,2'bx1} : dec_pc_set_op01 = 1'b1;  /* SOFT2,,BREAK */
                {8'h61,8'hb1,2'bx1} : dec_pc_set_op01 = 1'b1;  /* SOFT3,,BREAK */
                {8'h61,8'hc1,2'bx1} : dec_pc_set_op01 = 1'b1;  /* SOFT4,,BREAK */
                default : dec_pc_set_op01 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_pc_set_op12;
    reg    dec_pc_set_op12;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_pc_set_op12 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'hfd,8'hxx,2'bx0} : dec_pc_set_op12 = 1'b1;  /* CALL,,!addr16 */
                {8'hed,8'hxx,2'bx0} : dec_pc_set_op12 = 1'b1;  /* BR,,!addr16 */
                default : dec_pc_set_op12 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_pc_set_op123;
    reg    dec_pc_set_op123;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_pc_set_op123 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'hfc,8'hxx,2'bx0} : dec_pc_set_op123 = 1'b1;  /* CALL,,!!addr20 */
                {8'hec,8'hxx,2'bx0} : dec_pc_set_op123 = 1'b1;  /* BR,,!!addr20 */
                default : dec_pc_set_op123 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_pc_set_AX;
    reg    dec_pc_set_AX;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_pc_set_AX = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hca,2'bx0} : dec_pc_set_AX = 1'b1;  /* CALL,,AX */
                {8'h61,8'hcb,2'bx0} : dec_pc_set_AX = 1'b1;  /* BR,,AX */
                default : dec_pc_set_AX = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_pc_set_BC;
    reg    dec_pc_set_BC;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_pc_set_BC = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hda,2'bx0} : dec_pc_set_BC = 1'b1;  /* CALL,,BC */
                default : dec_pc_set_BC = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_pc_set_DE;
    reg    dec_pc_set_DE;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_pc_set_DE = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hea,2'bx0} : dec_pc_set_DE = 1'b1;  /* CALL,,DE */
                default : dec_pc_set_DE = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_pc_set_HL;
    reg    dec_pc_set_HL;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_pc_set_HL = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hfa,2'bx0} : dec_pc_set_HL = 1'b1;  /* CALL,,HL */
                default : dec_pc_set_HL = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_pc_set_pc1;
    reg    dec_pc_set_pc1;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_pc_set_pc1 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'hef,8'hxx,2'bx0} : dec_pc_set_pc1 = 1'b1;  /* BR,,$addr8 */
                {8'hdc,8'hxx,2'bx1} : dec_pc_set_pc1 = 1'b1;  /* BC,,$addr8 */
                {8'hde,8'hxx,2'bx1} : dec_pc_set_pc1 = 1'b1;  /* BNC,,$addr8 */
                {8'hdd,8'hxx,2'bx1} : dec_pc_set_pc1 = 1'b1;  /* BZ,,$addr8 */
                {8'hdf,8'hxx,2'bx1} : dec_pc_set_pc1 = 1'b1;  /* BNZ,,$addr8 */
                default : dec_pc_set_pc1 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_pc_set_pc2;
    reg    dec_pc_set_pc2;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_pc_set_pc2 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hc3,2'bx1} : dec_pc_set_pc2 = 1'b1;  /* BH,,$addr8 */
                {8'h61,8'hd3,2'bx1} : dec_pc_set_pc2 = 1'b1;  /* BNH,,$addr8 */
                {8'h31,8'h03,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BT,A.0,$addr8 */
                {8'h31,8'h13,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BT,A.1,$addr8 */
                {8'h31,8'h23,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BT,A.2,$addr8 */
                {8'h31,8'h33,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BT,A.3,$addr8 */
                {8'h31,8'h43,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BT,A.4,$addr8 */
                {8'h31,8'h53,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BT,A.5,$addr8 */
                {8'h31,8'h63,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BT,A.6,$addr8 */
                {8'h31,8'h73,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BT,A.7,$addr8 */
                {8'h31,8'h83,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BT,[HL].0,$addr8 */
                {8'h31,8'h93,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BT,[HL].1,$addr8 */
                {8'h31,8'ha3,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BT,[HL].2,$addr8 */
                {8'h31,8'hb3,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BT,[HL].3,$addr8 */
                {8'h31,8'hc3,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BT,[HL].4,$addr8 */
                {8'h31,8'hd3,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BT,[HL].5,$addr8 */
                {8'h31,8'he3,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BT,[HL].6,$addr8 */
                {8'h31,8'hf3,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BT,[HL].7,$addr8 */
                {8'h31,8'h05,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BF,A.0,$addr8 */
                {8'h31,8'h15,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BF,A.1,$addr8 */
                {8'h31,8'h25,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BF,A.2,$addr8 */
                {8'h31,8'h35,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BF,A.3,$addr8 */
                {8'h31,8'h45,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BF,A.4,$addr8 */
                {8'h31,8'h55,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BF,A.5,$addr8 */
                {8'h31,8'h65,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BF,A.6,$addr8 */
                {8'h31,8'h75,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BF,A.7,$addr8 */
                {8'h31,8'h85,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BF,[HL].0,$addr8 */
                {8'h31,8'h95,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BF,[HL].1,$addr8 */
                {8'h31,8'ha5,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BF,[HL].2,$addr8 */
                {8'h31,8'hb5,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BF,[HL].3,$addr8 */
                {8'h31,8'hc5,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BF,[HL].4,$addr8 */
                {8'h31,8'hd5,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BF,[HL].5,$addr8 */
                {8'h31,8'he5,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BF,[HL].6,$addr8 */
                {8'h31,8'hf5,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BF,[HL].7,$addr8 */
                {8'h31,8'h01,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BTCLR,A.0,$addr8 */
                {8'h31,8'h11,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BTCLR,A.1,$addr8 */
                {8'h31,8'h21,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BTCLR,A.2,$addr8 */
                {8'h31,8'h31,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BTCLR,A.3,$addr8 */
                {8'h31,8'h41,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BTCLR,A.4,$addr8 */
                {8'h31,8'h51,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BTCLR,A.5,$addr8 */
                {8'h31,8'h61,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BTCLR,A.6,$addr8 */
                {8'h31,8'h71,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BTCLR,A.7,$addr8 */
                {8'h31,8'h81,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BTCLR,[HL].0,$addr8 */
                {8'h31,8'h91,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BTCLR,[HL].1,$addr8 */
                {8'h31,8'ha1,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BTCLR,[HL].2,$addr8 */
                {8'h31,8'hb1,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BTCLR,[HL].3,$addr8 */
                {8'h31,8'hc1,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BTCLR,[HL].4,$addr8 */
                {8'h31,8'hd1,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BTCLR,[HL].5,$addr8 */
                {8'h31,8'he1,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BTCLR,[HL].6,$addr8 */
                {8'h31,8'hf1,2'b10} : dec_pc_set_pc2 = 1'b1;  /* BTCLR,[HL].7,$addr8 */
                default : dec_pc_set_pc2 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_pc_set_pc3;
    reg    dec_pc_set_pc3;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_pc_set_pc3 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h31,8'h02,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BT,saddr.0,$addr8 */
                {8'h31,8'h12,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BT,saddr.1,$addr8 */
                {8'h31,8'h22,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BT,saddr.2,$addr8 */
                {8'h31,8'h32,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BT,saddr.3,$addr8 */
                {8'h31,8'h42,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BT,saddr.4,$addr8 */
                {8'h31,8'h52,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BT,saddr.5,$addr8 */
                {8'h31,8'h62,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BT,saddr.6,$addr8 */
                {8'h31,8'h72,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BT,saddr.7,$addr8 */
                {8'h31,8'h82,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BT,sfr.0,$addr8 */
                {8'h31,8'h92,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BT,sfr.1,$addr8 */
                {8'h31,8'ha2,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BT,sfr.2,$addr8 */
                {8'h31,8'hb2,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BT,sfr.3,$addr8 */
                {8'h31,8'hc2,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BT,sfr.4,$addr8 */
                {8'h31,8'hd2,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BT,sfr.5,$addr8 */
                {8'h31,8'he2,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BT,sfr.6,$addr8 */
                {8'h31,8'hf2,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BT,sfr.7,$addr8 */
                {8'h31,8'h04,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BF,saddr.0,$addr8 */
                {8'h31,8'h14,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BF,saddr.1,$addr8 */
                {8'h31,8'h24,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BF,saddr.2,$addr8 */
                {8'h31,8'h34,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BF,saddr.3,$addr8 */
                {8'h31,8'h44,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BF,saddr.4,$addr8 */
                {8'h31,8'h54,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BF,saddr.5,$addr8 */
                {8'h31,8'h64,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BF,saddr.6,$addr8 */
                {8'h31,8'h74,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BF,saddr.7,$addr8 */
                {8'h31,8'h84,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BF,sfr.0,$addr8 */
                {8'h31,8'h94,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BF,sfr.1,$addr8 */
                {8'h31,8'ha4,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BF,sfr.2,$addr8 */
                {8'h31,8'hb4,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BF,sfr.3,$addr8 */
                {8'h31,8'hc4,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BF,sfr.4,$addr8 */
                {8'h31,8'hd4,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BF,sfr.5,$addr8 */
                {8'h31,8'he4,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BF,sfr.6,$addr8 */
                {8'h31,8'hf4,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BF,sfr.7,$addr8 */
                {8'h31,8'h00,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BTCLR,saddr.0,$addr8 */
                {8'h31,8'h10,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BTCLR,saddr.1,$addr8 */
                {8'h31,8'h20,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BTCLR,saddr.2,$addr8 */
                {8'h31,8'h30,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BTCLR,saddr.3,$addr8 */
                {8'h31,8'h40,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BTCLR,saddr.4,$addr8 */
                {8'h31,8'h50,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BTCLR,saddr.5,$addr8 */
                {8'h31,8'h60,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BTCLR,saddr.6,$addr8 */
                {8'h31,8'h70,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BTCLR,saddr.7,$addr8 */
                {8'h31,8'h80,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BTCLR,sfr.0,$addr8 */
                {8'h31,8'h90,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BTCLR,sfr.1,$addr8 */
                {8'h31,8'ha0,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BTCLR,sfr.2,$addr8 */
                {8'h31,8'hb0,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BTCLR,sfr.3,$addr8 */
                {8'h31,8'hc0,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BTCLR,sfr.4,$addr8 */
                {8'h31,8'hd0,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BTCLR,sfr.5,$addr8 */
                {8'h31,8'he0,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BTCLR,sfr.6,$addr8 */
                {8'h31,8'hf0,2'b10} : dec_pc_set_pc3 = 1'b1;  /* BTCLR,sfr.7,$addr8 */
                default : dec_pc_set_pc3 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_pc_set_pc12;
    reg    dec_pc_set_pc12;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_pc_set_pc12 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'hfe,8'hxx,2'bx0} : dec_pc_set_pc12 = 1'b1;  /* CALL,,$!addr16 */
                {8'hee,8'hxx,2'bx0} : dec_pc_set_pc12 = 1'b1;  /* BR,,$!addr16 */
                default : dec_pc_set_pc12 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_pc_set_calt;
    reg    dec_pc_set_calt;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_pc_set_calt = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'h84,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[0080h] */
                {8'h61,8'h94,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[0082h] */
                {8'h61,8'ha4,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[0084h] */
                {8'h61,8'hb4,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[0086h] */
                {8'h61,8'hc4,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[0088h] */
                {8'h61,8'hd4,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[008Ah] */
                {8'h61,8'he4,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[008Ch] */
                {8'h61,8'hf4,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[008Eh] */
                {8'h61,8'h85,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[0090h] */
                {8'h61,8'h95,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[0092h] */
                {8'h61,8'ha5,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[0094h] */
                {8'h61,8'hb5,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[0096h] */
                {8'h61,8'hc5,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[0098h] */
                {8'h61,8'hd5,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[009Ah] */
                {8'h61,8'he5,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[009Ch] */
                {8'h61,8'hf5,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[009Eh] */
                {8'h61,8'h86,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[00A0h] */
                {8'h61,8'h96,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[00A2h] */
                {8'h61,8'ha6,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[00A4h] */
                {8'h61,8'hb6,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[00A6h] */
                {8'h61,8'hc6,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[00A8h] */
                {8'h61,8'hd6,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[00AAh] */
                {8'h61,8'he6,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[00ACh] */
                {8'h61,8'hf6,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[00AEh] */
                {8'h61,8'h87,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[00B0h] */
                {8'h61,8'h97,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[00B2h] */
                {8'h61,8'ha7,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[00B4h] */
                {8'h61,8'hb7,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[00B6h] */
                {8'h61,8'hc7,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[00B8h] */
                {8'h61,8'hd7,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[00BAh] */
                {8'h61,8'he7,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[00BCh] */
                {8'h61,8'hf7,2'bx0} : dec_pc_set_calt = 1'b1;  /* CALLT,,[00BEh] */
                default : dec_pc_set_calt = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_pc_set_vec;
    reg    dec_pc_set_vec;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(decout_mask == 1'b1) begin
//            dec_pc_set_vec = 1'b0;
//        end else if(rstvec == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1) begin
            dec_pc_set_vec = 1'b0;
        end else if(ivack == 1'b1) begin
            casex ({stage_adr})  
                {2'b01} : dec_pc_set_vec = 1'b1;  /* Interrupt */
                default : dec_pc_set_vec = 1'b0;
            endcase
        end else if(skpack == 1'b1) begin
            dec_pc_set_vec = 1'b0;
        end else begin
            dec_pc_set_vec = 1'b0;
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_pc_set_brk;
    reg    dec_pc_set_brk;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_pc_set_brk = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hcc,2'bx0} : dec_pc_set_brk = 1'b1;  /* BRK,, */
                default : dec_pc_set_brk = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_pc_set_ret;
    reg    dec_pc_set_ret;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_pc_set_ret = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'hd7,8'hxx,2'b11} : dec_pc_set_ret = 1'b1;  /* RET,, */
                {8'h61,8'hec,2'b11} : dec_pc_set_ret = 1'b1;  /* RETB,, */
                {8'h61,8'hfc,2'b11} : dec_pc_set_ret = 1'b1;  /* RETI,, */
                default : dec_pc_set_ret = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_pc_set_dbg;
    reg    dec_pc_set_dbg;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_pc_set_dbg = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'hff,8'hxx,2'bx0} : dec_pc_set_dbg = 1'b1;  /* SOFT,,BREAK */
                {8'h61,8'ha1,2'bx0} : dec_pc_set_dbg = 1'b1;  /* SOFT2,,BREAK */
                {8'h61,8'hb1,2'bx0} : dec_pc_set_dbg = 1'b1;  /* SOFT3,,BREAK */
                {8'h61,8'hc1,2'bx0} : dec_pc_set_dbg = 1'b1;  /* SOFT4,,BREAK */
                default : dec_pc_set_dbg = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_stage_cut_brtf;
    reg    dec_stage_cut_brtf;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_stage_cut_brtf = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h31,8'h02,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,saddr.0,$addr8 */
                {8'h31,8'h12,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,saddr.1,$addr8 */
                {8'h31,8'h22,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,saddr.2,$addr8 */
                {8'h31,8'h32,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,saddr.3,$addr8 */
                {8'h31,8'h42,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,saddr.4,$addr8 */
                {8'h31,8'h52,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,saddr.5,$addr8 */
                {8'h31,8'h62,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,saddr.6,$addr8 */
                {8'h31,8'h72,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,saddr.7,$addr8 */
                {8'h31,8'h82,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,sfr.0,$addr8 */
                {8'h31,8'h92,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,sfr.1,$addr8 */
                {8'h31,8'ha2,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,sfr.2,$addr8 */
                {8'h31,8'hb2,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,sfr.3,$addr8 */
                {8'h31,8'hc2,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,sfr.4,$addr8 */
                {8'h31,8'hd2,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,sfr.5,$addr8 */
                {8'h31,8'he2,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,sfr.6,$addr8 */
                {8'h31,8'hf2,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,sfr.7,$addr8 */
                {8'h31,8'h03,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,A.0,$addr8 */
                {8'h31,8'h13,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,A.1,$addr8 */
                {8'h31,8'h23,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,A.2,$addr8 */
                {8'h31,8'h33,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,A.3,$addr8 */
                {8'h31,8'h43,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,A.4,$addr8 */
                {8'h31,8'h53,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,A.5,$addr8 */
                {8'h31,8'h63,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,A.6,$addr8 */
                {8'h31,8'h73,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,A.7,$addr8 */
                {8'h31,8'h83,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,[HL].0,$addr8 */
                {8'h31,8'h93,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,[HL].1,$addr8 */
                {8'h31,8'ha3,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,[HL].2,$addr8 */
                {8'h31,8'hb3,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,[HL].3,$addr8 */
                {8'h31,8'hc3,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,[HL].4,$addr8 */
                {8'h31,8'hd3,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,[HL].5,$addr8 */
                {8'h31,8'he3,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,[HL].6,$addr8 */
                {8'h31,8'hf3,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BT,[HL].7,$addr8 */
                {8'h31,8'h04,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,saddr.0,$addr8 */
                {8'h31,8'h14,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,saddr.1,$addr8 */
                {8'h31,8'h24,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,saddr.2,$addr8 */
                {8'h31,8'h34,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,saddr.3,$addr8 */
                {8'h31,8'h44,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,saddr.4,$addr8 */
                {8'h31,8'h54,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,saddr.5,$addr8 */
                {8'h31,8'h64,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,saddr.6,$addr8 */
                {8'h31,8'h74,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,saddr.7,$addr8 */
                {8'h31,8'h84,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,sfr.0,$addr8 */
                {8'h31,8'h94,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,sfr.1,$addr8 */
                {8'h31,8'ha4,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,sfr.2,$addr8 */
                {8'h31,8'hb4,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,sfr.3,$addr8 */
                {8'h31,8'hc4,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,sfr.4,$addr8 */
                {8'h31,8'hd4,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,sfr.5,$addr8 */
                {8'h31,8'he4,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,sfr.6,$addr8 */
                {8'h31,8'hf4,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,sfr.7,$addr8 */
                {8'h31,8'h05,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,A.0,$addr8 */
                {8'h31,8'h15,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,A.1,$addr8 */
                {8'h31,8'h25,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,A.2,$addr8 */
                {8'h31,8'h35,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,A.3,$addr8 */
                {8'h31,8'h45,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,A.4,$addr8 */
                {8'h31,8'h55,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,A.5,$addr8 */
                {8'h31,8'h65,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,A.6,$addr8 */
                {8'h31,8'h75,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,A.7,$addr8 */
                {8'h31,8'h85,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,[HL].0,$addr8 */
                {8'h31,8'h95,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,[HL].1,$addr8 */
                {8'h31,8'ha5,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,[HL].2,$addr8 */
                {8'h31,8'hb5,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,[HL].3,$addr8 */
                {8'h31,8'hc5,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,[HL].4,$addr8 */
                {8'h31,8'hd5,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,[HL].5,$addr8 */
                {8'h31,8'he5,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,[HL].6,$addr8 */
                {8'h31,8'hf5,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BF,[HL].7,$addr8 */
                {8'h31,8'h00,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,saddr.0,$addr8 */
                {8'h31,8'h10,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,saddr.1,$addr8 */
                {8'h31,8'h20,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,saddr.2,$addr8 */
                {8'h31,8'h30,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,saddr.3,$addr8 */
                {8'h31,8'h40,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,saddr.4,$addr8 */
                {8'h31,8'h50,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,saddr.5,$addr8 */
                {8'h31,8'h60,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,saddr.6,$addr8 */
                {8'h31,8'h70,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,saddr.7,$addr8 */
                {8'h31,8'h80,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,sfr.0,$addr8 */
                {8'h31,8'h90,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,sfr.1,$addr8 */
                {8'h31,8'ha0,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,sfr.2,$addr8 */
                {8'h31,8'hb0,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,sfr.3,$addr8 */
                {8'h31,8'hc0,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,sfr.4,$addr8 */
                {8'h31,8'hd0,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,sfr.5,$addr8 */
                {8'h31,8'he0,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,sfr.6,$addr8 */
                {8'h31,8'hf0,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,sfr.7,$addr8 */
                {8'h31,8'h01,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,A.0,$addr8 */
                {8'h31,8'h11,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,A.1,$addr8 */
                {8'h31,8'h21,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,A.2,$addr8 */
                {8'h31,8'h31,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,A.3,$addr8 */
                {8'h31,8'h41,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,A.4,$addr8 */
                {8'h31,8'h51,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,A.5,$addr8 */
                {8'h31,8'h61,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,A.6,$addr8 */
                {8'h31,8'h71,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,A.7,$addr8 */
                {8'h31,8'h81,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,[HL].0,$addr8 */
                {8'h31,8'h91,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,[HL].1,$addr8 */
                {8'h31,8'ha1,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,[HL].2,$addr8 */
                {8'h31,8'hb1,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,[HL].3,$addr8 */
                {8'h31,8'hc1,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,[HL].4,$addr8 */
                {8'h31,8'hd1,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,[HL].5,$addr8 */
                {8'h31,8'he1,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,[HL].6,$addr8 */
                {8'h31,8'hf1,2'b01} : dec_stage_cut_brtf = 1'b1;  /* BTCLR,[HL].7,$addr8 */
                default : dec_stage_cut_brtf = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_stage_cut_ifbr;
    reg    dec_stage_cut_ifbr;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_stage_cut_ifbr = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'hdc,8'hxx,2'bx0} : dec_stage_cut_ifbr = 1'b1;  /* BC,,$addr8 */
                {8'hde,8'hxx,2'bx0} : dec_stage_cut_ifbr = 1'b1;  /* BNC,,$addr8 */
                {8'hdd,8'hxx,2'bx0} : dec_stage_cut_ifbr = 1'b1;  /* BZ,,$addr8 */
                {8'hdf,8'hxx,2'bx0} : dec_stage_cut_ifbr = 1'b1;  /* BNZ,,$addr8 */
                {8'h61,8'hc3,2'bx0} : dec_stage_cut_ifbr = 1'b1;  /* BH,,$addr8 */
                {8'h61,8'hd3,2'bx0} : dec_stage_cut_ifbr = 1'b1;  /* BNH,,$addr8 */
                default : dec_stage_cut_ifbr = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ifbr_not;
    reg    dec_ifbr_not;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_ifbr_not = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'hde,8'hxx,2'bx0} : dec_ifbr_not = 1'b1;  /* BNC,,$addr8 */
                {8'hdf,8'hxx,2'bx0} : dec_ifbr_not = 1'b1;  /* BNZ,,$addr8 */
                {8'h61,8'hd3,2'bx0} : dec_ifbr_not = 1'b1;  /* BNH,,$addr8 */
                default : dec_ifbr_not = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ifbr_zero;
    reg    dec_ifbr_zero;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_ifbr_zero = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'hdd,8'hxx,2'bx0} : dec_ifbr_zero = 1'b1;  /* BZ,,$addr8 */
                {8'hdf,8'hxx,2'bx0} : dec_ifbr_zero = 1'b1;  /* BNZ,,$addr8 */
                default : dec_ifbr_zero = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_ifbr_ht;
    reg    dec_ifbr_ht;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_ifbr_ht = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hc3,2'bx0} : dec_ifbr_ht = 1'b1;  /* BH,,$addr8 */
                {8'h61,8'hd3,2'bx0} : dec_ifbr_ht = 1'b1;  /* BNH,,$addr8 */
                default : dec_ifbr_ht = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_mem_stage_op2;
    reg    dec_mem_stage_op2;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_mem_stage_op2 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1})  
                {8'hcd,8'hxx} : dec_mem_stage_op2 = 1'b1;  /* MOV,saddr,#byte */
                {8'hce,8'hxx} : dec_mem_stage_op2 = 1'b1;  /* MOV,sfr,#byte */
                {8'hca,8'hxx} : dec_mem_stage_op2 = 1'b1;  /* MOV,[DE+byte],#byte */
                {8'hcc,8'hxx} : dec_mem_stage_op2 = 1'b1;  /* MOV,[HL+byte],#byte */
                {8'hc8,8'hxx} : dec_mem_stage_op2 = 1'b1;  /* MOV,[SP+byte],#byte */
                {8'h0a,8'hxx} : dec_mem_stage_op2 = 1'b1;  /* ADD,saddr,#byte */
                {8'h1a,8'hxx} : dec_mem_stage_op2 = 1'b1;  /* ADDC,saddr,#byte */
                {8'h2a,8'hxx} : dec_mem_stage_op2 = 1'b1;  /* SUB,saddr,#byte */
                {8'h3a,8'hxx} : dec_mem_stage_op2 = 1'b1;  /* SUBC,saddr,#byte */
                {8'h5a,8'hxx} : dec_mem_stage_op2 = 1'b1;  /* AND,saddr,#byte */
                {8'h6a,8'hxx} : dec_mem_stage_op2 = 1'b1;  /* OR,saddr,#byte */
                {8'h7a,8'hxx} : dec_mem_stage_op2 = 1'b1;  /* XOR,saddr,#byte */
                {8'h4a,8'hxx} : dec_mem_stage_op2 = 1'b1;  /* CMP,saddr,#byte */
                default : dec_mem_stage_op2 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_mem_stage_op3;
    reg    dec_mem_stage_op3;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_mem_stage_op3 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1})  
                {8'hcf,8'hxx} : dec_mem_stage_op3 = 1'b1;  /* MOV,!addr16,#byte */
                {8'h19,8'hxx} : dec_mem_stage_op3 = 1'b1;  /* MOV,word[B],#byte */
                {8'h38,8'hxx} : dec_mem_stage_op3 = 1'b1;  /* MOV,word[C],#byte */
                {8'h39,8'hxx} : dec_mem_stage_op3 = 1'b1;  /* MOV,word[BC],#byte */
                {8'h40,8'hxx} : dec_mem_stage_op3 = 1'b1;  /* CMP,!addr16,#byte */
                default : dec_mem_stage_op3 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_mem_stage_op23;
    reg    dec_mem_stage_op23;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_mem_stage_op23 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1})  
                {8'hc9,8'hxx} : dec_mem_stage_op23 = 1'b1;  /* MOVW,saddrp,#word */
                {8'hcb,8'hxx} : dec_mem_stage_op23 = 1'b1;  /* MOVW,sfrp,#word */
                default : dec_mem_stage_op23 = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_set_buf_retadr;
    reg    dec_set_buf_retadr;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_set_buf_retadr = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hca,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALL,,AX */
                {8'h61,8'hda,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALL,,BC */
                {8'h61,8'hea,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALL,,DE */
                {8'h61,8'hfa,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALL,,HL */
                {8'hfe,8'hxx,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALL,,$!addr16 */
                {8'hfd,8'hxx,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALL,,!addr16 */
                {8'hfc,8'hxx,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALL,,!!addr20 */
                {8'h61,8'h84,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[0080h] */
                {8'h61,8'h94,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[0082h] */
                {8'h61,8'ha4,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[0084h] */
                {8'h61,8'hb4,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[0086h] */
                {8'h61,8'hc4,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[0088h] */
                {8'h61,8'hd4,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[008Ah] */
                {8'h61,8'he4,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[008Ch] */
                {8'h61,8'hf4,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[008Eh] */
                {8'h61,8'h85,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[0090h] */
                {8'h61,8'h95,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[0092h] */
                {8'h61,8'ha5,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[0094h] */
                {8'h61,8'hb5,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[0096h] */
                {8'h61,8'hc5,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[0098h] */
                {8'h61,8'hd5,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[009Ah] */
                {8'h61,8'he5,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[009Ch] */
                {8'h61,8'hf5,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[009Eh] */
                {8'h61,8'h86,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[00A0h] */
                {8'h61,8'h96,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[00A2h] */
                {8'h61,8'ha6,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[00A4h] */
                {8'h61,8'hb6,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[00A6h] */
                {8'h61,8'hc6,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[00A8h] */
                {8'h61,8'hd6,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[00AAh] */
                {8'h61,8'he6,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[00ACh] */
                {8'h61,8'hf6,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[00AEh] */
                {8'h61,8'h87,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[00B0h] */
                {8'h61,8'h97,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[00B2h] */
                {8'h61,8'ha7,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[00B4h] */
                {8'h61,8'hb7,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[00B6h] */
                {8'h61,8'hc7,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[00B8h] */
                {8'h61,8'hd7,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[00BAh] */
                {8'h61,8'he7,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[00BCh] */
                {8'h61,8'hf7,2'bx0} : dec_set_buf_retadr = 1'b1;  /* CALLT,,[00BEh] */
                {8'h61,8'hcc,2'bx0} : dec_set_buf_retadr = 1'b1;  /* BRK,, */
                {8'hff,8'hxx,2'bx0} : dec_set_buf_retadr = 1'b1;  /* SOFT,,BREAK */
                {8'h61,8'ha1,2'bx0} : dec_set_buf_retadr = 1'b1;  /* SOFT2,,BREAK */
                {8'h61,8'hb1,2'bx0} : dec_set_buf_retadr = 1'b1;  /* SOFT3,,BREAK */
                {8'h61,8'hc1,2'bx0} : dec_set_buf_retadr = 1'b1;  /* SOFT4,,BREAK */
                default : dec_set_buf_retadr = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_set_buf_intr;
    reg    dec_set_buf_intr;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(decout_mask == 1'b1) begin
//            dec_set_buf_intr = 1'b0;
//        end else if(rstvec == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1) begin
            dec_set_buf_intr = 1'b0;
        end else if(ivack == 1'b1) begin
            casex ({stage_adr}) 
                 {2'b00} : dec_set_buf_intr = 1'b1;  /* Interrupt */
                default : dec_set_buf_intr = 1'b0;
            endcase
        end else if(skpack == 1'b1) begin
            dec_set_buf_intr = 1'b0;
        end else begin
            dec_set_buf_intr = 1'b0;
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_skc;
    reg    dec_skc;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_skc = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr}) 
                 {8'h61,8'hc8,2'bxx} : dec_skc = 1'b1;  /* SKC,, */
                default : dec_skc = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_sknc;
    reg    dec_sknc;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_sknc = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr}) 
                 {8'h61,8'hd8,2'bxx} : dec_sknc = 1'b1;  /* SKNC,, */
                default : dec_sknc = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_skz;
    reg    dec_skz;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_skz = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr}) 
                 {8'h61,8'he8,2'bxx} : dec_skz = 1'b1;  /* SKZ,, */
                default : dec_skz = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_sknz;
    reg    dec_sknz;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_sknz = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr}) 
                 {8'h61,8'hf8,2'bxx} : dec_sknz = 1'b1;  /* SKNZ,, */
                default : dec_sknz = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_skh;
    reg    dec_skh;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_skh = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr}) 
                 {8'h61,8'he3,2'bxx} : dec_skh = 1'b1;  /* SKH,, */
                default : dec_skh = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_sknh;
    reg    dec_sknh;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_sknh = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr}) 
                 {8'h61,8'hf3,2'bxx} : dec_sknh = 1'b1;  /* SKNH,, */
                default : dec_sknh = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_prefix;
    reg    dec_prefix;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_prefix = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h11,8'hxx,2'bxx} : dec_prefix = 1'b1;  /* PREFIX,, */
                default : dec_prefix = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_halt;
    reg    dec_halt;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_halt = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hed,2'b01} : dec_halt = 1'b1;  /* HALT,, */
                default : dec_halt = 1'b0;
            endcase
        end
    end

/*------------------------------------------------------------------------------*/
/* Ver2.0  									*/
/*�����ǥ��������Ϥ�decout_mask�ǥޥ������롣					*/
/*------------------------------------------------------------------------------*/

    output dec_stop;
    reg    dec_stop;
//    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack or decout_mask) begin
//        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1 || decout_mask == 1'b1) begin
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_stop = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hfd,2'b01} : dec_stop = 1'b1;  /* STOP,, */
                default : dec_stop = 1'b0;
            endcase
        end
    end
    output dec_movs;
    reg    dec_movs, dec_movs_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_movs_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hce,2'bxx} : dec_movs_adrstage = 1'b1;  /* MOVS,[HL+byte],X */
                default : dec_movs_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_movs <= 1'b0;
        else if(cpuen) dec_movs <= dec_movs_adrstage;
    end
    output dec_cmps;
    reg    dec_cmps, dec_cmps_adrstage;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_cmps_adrstage = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'hde,2'bxx} : dec_cmps_adrstage = 1'b1;  /* CMPS,X,[HL+byte] */
                default : dec_cmps_adrstage = 1'b0;
            endcase
        end
    end
    //synopsys async_set_reset "resb"
    always @(posedge baseck or negedge resb) begin
        if (!resb) dec_cmps <= 1'b0;
        else if(cpuen) dec_cmps <= dec_cmps_adrstage;
    end

// for EVA
    output dec_alt1;
    reg    dec_alt1;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_alt1 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'h81,2'bxx} : dec_alt1 = 1'b1;  /* ALT1,, */
                default : dec_alt1 = 1'b0;
            endcase
        end
    end
    output dec_alt2;
    reg    dec_alt2;
    always @(ID_stage0 or ID_stage1 or stage_adr or ivack or rstvec or skpack) begin
        if(rstvec == 1'b1 || ivack == 1'b1 || skpack == 1'b1) begin
            dec_alt2 = 1'b0;
        end else begin
            casex ({ID_stage0,ID_stage1,stage_adr})  
                {8'h61,8'h91,2'bxx} : dec_alt2 = 1'b1;  /* ALT2,, */
                default : dec_alt2 = 1'b0;
            endcase
        end
    end
//

endmodule

/*--------------------------------------------------------------------------------------*/
/* Ver2.0  										*/
/*  �ǥ������ν��Ϥ�ޥ�������ǥ��쥤�ǻҡ�						*/
//��TBDLY2X2�Ϣ�1.8502ns, ��1.5337ns���ǥ��������ٱ䤬��7ns�Ǥ��뤿�ᡢ���Ĥ���Ѥ��롣	*/
//���ٱ��ͤϥǥ������ν����ٱ��ǥ��쥤�ǻҤȤʤ������				*/
//���������ٱ�򥪡��С����Ƥ���ή������������Τ��ᡢ9�����٤Υǥ��������Ϥ򥫥С�	*/
//������Ф褯���ü��������դ��ʤ���Dont tuch�����Ȥ��롣				*/
//�������ٱ��SLFLASH�η�ϩ�ǥ��ԡ��ɥͥå��ѥ��Ȥʤ뤿�ᡢ�ǹ�®�������(DECDYCUT=1)��	*/
//�����Ϥ��β�ϩ��ư���ʤ��褦�ˤ��롣							*/
//���ץ������Ѥ�ä��ݤϾ嵭���򸵤�Ĵ�����뤳�ȡ�					*/
/*--------------------------------------------------------------------------------------*/
/* Ver3.0 �ǥ��쥤�ˤ��ҥ��ɻ߲�ϩ���к���ľ��(CPUv1.5���������᤹)		*/
/*------------------------------------------------------------------------------*/
//module QLK0RCPUEVA0V3_DEC_DLY(out, in);
//	input in;
//	output out;
// // for EVA
// //	wire net1, net2, net3, net4;
// //	TBDLY2X2 dly1 ( .N01(net1), .H01(in)   );
// //	TBDLY2X2 dly2 ( .N01(net2), .H01(net1) );
// //	TBDLY2X2 dly3 ( .N01(net3), .H01(net2) );
// //	TBDLY2X2 dly4 ( .N01(net4), .H01(net3) );
// //	TBDLY2X2 dly5 ( .N01(out),  .H01(net4) );
//
// // for EVA
//        assign out = in ;
//
//
//endmodule


module da_ICE(da_data,FMAIN_FCLK,FCLK);  
   input [1:0] da_data;
   output 	   FMAIN_FCLK;
   output      FCLK;
   
endmodule // da_ICE

module m1767_ff3(RESB,O,VIMDS1,VIMDS0);
   input RESB;
   output O;
   input  VIMDS1,VIMDS0;
   
   assign RESB = O;   
endmodule // 1767_ff3

/****************************************************************/
/* Date		: 2007/10/12					*/
/* Revision	: 1.00						*/
/* Designer	: T.Tsunoda					*/
/****************************************************************/

module	icescon (
		TIIDER, ICEMSKCKSMER, CKSMER, PSEUDOCKSMER,
		CSPDTFLP,
		ICEIFA31, ICEIFA30, ICEIFA29, ICEIFA28, ICEIFA27, ICEIFA26, ICEIFA25, ICEIFA24,
		ICEIFA23, ICEIFA22, ICEIFA21, ICEIFA20, ICEIFA19, ICEIFA18, ICEIFA17, ICEIFA16,
		ICEIFA15, ICEIFA14, ICEIFA13, ICEIFA12, ICEIFA11, ICEIFA10, ICEIFA9,  ICEIFA8,
		ICEIFA7,  ICEIFA6,  ICEIFA5,  ICEIFA4,  ICEIFA3,  ICEIFA2,  ICEIFA1,  ICEIFA0,
		ICEDI31, ICEDI30, ICEDI29, ICEDI28, ICEDI27, ICEDI26, ICEDI25, ICEDI24,
		ICEDI23, ICEDI22, ICEDI21, ICEDI20, ICEDI19, ICEDI18, ICEDI17, ICEDI16,
		ICEDI15, ICEDI14, ICEDI13, ICEDI12, ICEDI11, ICEDI10, ICEDI9,  ICEDI8,
		ICEDI7,  ICEDI6,  ICEDI5,  ICEDI4,  ICEDI3,  ICEDI2,  ICEDI1,  ICEDI0,
		ICEWR, FCLKRT, SYSRSOUTB,
		ICEDOP31, ICEDOP30, ICEDOP29, ICEDOP28, ICEDOP27, ICEDOP26, ICEDOP25, ICEDOP24,
		ICEDOP23, ICEDOP22, ICEDOP21, ICEDOP20, ICEDOP19, ICEDOP18, ICEDOP17, ICEDOP16,
		ICEDOP15, ICEDOP14, ICEDOP13, ICEDOP12, ICEDOP11, ICEDOP10, ICEDOP9,  ICEDOP8,
		ICEDOP7,  ICEDOP6,  ICEDOP5,  ICEDOP4,  ICEDOP3,  ICEDOP2,  ICEDOP1,  ICEDOP0,
		ICECKSMER, CSPDTFLG
		);

	input	TIIDER;					// mode��˥��к�
	input	ICEMSKCKSMER, CKSMER, PSEUDOCKSMER;	// cib sec
	input	CSPDTFLP;
	input	ICEIFA31, ICEIFA30, ICEIFA29, ICEIFA28, ICEIFA27, ICEIFA26, ICEIFA25, ICEIFA24,
		ICEIFA23, ICEIFA22, ICEIFA21, ICEIFA20, ICEIFA19, ICEIFA18, ICEIFA17, ICEIFA16,
		ICEIFA15, ICEIFA14, ICEIFA13, ICEIFA12, ICEIFA11, ICEIFA10, ICEIFA9,  ICEIFA8,
		ICEIFA7,  ICEIFA6,  ICEIFA5,  ICEIFA4,  ICEIFA3,  ICEIFA2,  ICEIFA1,  ICEIFA0;
	input	ICEDI31, ICEDI30, ICEDI29, ICEDI28, ICEDI27, ICEDI26, ICEDI25, ICEDI24,
		ICEDI23, ICEDI22, ICEDI21, ICEDI20, ICEDI19, ICEDI18, ICEDI17, ICEDI16,
		ICEDI15, ICEDI14, ICEDI13, ICEDI12, ICEDI11, ICEDI10, ICEDI9,  ICEDI8,
		ICEDI7,  ICEDI6,  ICEDI5,  ICEDI4,  ICEDI3,  ICEDI2,  ICEDI1,  ICEDI0;
	input	ICEWR, FCLKRT, SYSRSOUTB;
	output	ICECKSMER;
	output	CSPDTFLG;
	output	ICEDOP31, ICEDOP30, ICEDOP29, ICEDOP28, ICEDOP27, ICEDOP26, ICEDOP25, ICEDOP24,
		ICEDOP23, ICEDOP22, ICEDOP21, ICEDOP20, ICEDOP19, ICEDOP18, ICEDOP17, ICEDOP16,
		ICEDOP15, ICEDOP14, ICEDOP13, ICEDOP12, ICEDOP11, ICEDOP10, ICEDOP9,  ICEDOP8,
		ICEDOP7,  ICEDOP6,  ICEDOP5,  ICEDOP4,  ICEDOP3,  ICEDOP2,  ICEDOP1,  ICEDOP0;


	wire [31:0] icedi, icedo;
	assign	ICECKSMER = PSEUDOCKSMER | (ICEMSKCKSMER & CKSMER);

	wire	dfdiffcs = {
			ICEIFA31, ICEIFA30, ICEIFA29, ICEIFA28, ICEIFA27, ICEIFA26,
			ICEIFA25, ICEIFA24, ICEIFA23, ICEIFA22, ICEIFA21, ICEIFA20,
			ICEIFA19, ICEIFA18, ICEIFA17, ICEIFA16, ICEIFA15, ICEIFA14,
			ICEIFA13, ICEIFA12, ICEIFA11, ICEIFA10, ICEIFA9, ICEIFA8,
			ICEIFA7, ICEIFA6, ICEIFA5, ICEIFA4, ICEIFA3, ICEIFA2, 2'b00
		} == 32'h0400_0000;

	assign	icedi = {
			ICEDI31, ICEDI30, ICEDI29, ICEDI28, ICEDI27, ICEDI26,
			ICEDI25, ICEDI24, ICEDI23, ICEDI22, ICEDI21, ICEDI20,
			ICEDI19, ICEDI18, ICEDI17, ICEDI16, ICEDI15, ICEDI14,
			ICEDI13, ICEDI12, ICEDI11, ICEDI10, ICEDI9, ICEDI8,
			ICEDI7, ICEDI6, ICEDI5, ICEDI4, ICEDI3, ICEDI2,
			ICEDI1, ICEDI0
		};

	reg [31:0] dfdiffp2;
	always @(negedge ICEWR or negedge SYSRSOUTB) begin
		if (!SYSRSOUTB)		dfdiffp2 <= 32'h0;
		else if (dfdiffcs)	dfdiffp2 <= icedi;
	end
	reg [31:0] dfdiffp1;
	always @(posedge FCLKRT or negedge SYSRSOUTB) begin
		if (!SYSRSOUTB)	dfdiffp1 <= 32'h0;
		else		dfdiffp1 <= dfdiffp2;
	end
	reg [31:0] dfdiff;
	always @(posedge FCLKRT or negedge SYSRSOUTB) begin
		if (!SYSRSOUTB) dfdiff <= 32'h0;
		else		dfdiff <= dfdiffp1;
	end

	assign	CSPDTFLG = (dfdiff == 32'hffae_6832) ? CSPDTFLP : 1'b0;

	assign	icedo = dfdiffcs ? dfdiff : 32'h0;
	assign	{ICEDOP31, ICEDOP30, ICEDOP29, ICEDOP28, ICEDOP27, ICEDOP26, ICEDOP25, ICEDOP24,
		 ICEDOP23, ICEDOP22, ICEDOP21, ICEDOP20, ICEDOP19, ICEDOP18, ICEDOP17, ICEDOP16,
		 ICEDOP15, ICEDOP14, ICEDOP13, ICEDOP12, ICEDOP11, ICEDOP10, ICEDOP9, ICEDOP8,
		 ICEDOP7, ICEDOP6, ICEDOP5, ICEDOP4, ICEDOP3, ICEDOP2, ICEDOP1, ICEDOP0} = icedo;

endmodule

module svmodif(SVSTOP,SVSTOPICE);
   input SVSTOP;
   output SVSTOPICE;
   assign SVSTOPICE = SVSTOP;
endmodule
// ============================================================================================================	*/
/* K0R IECUBE ORBUS												*/
/* V100												tsunoda		*/
/* $Id: orbus-SS3rd.v,v 1.2 2010-02-01 02:59:25 snisimu Exp $							*/
/* ============================================================================================================	*/
module ORBUS (
	MDR_RAM15, MDR_RAM14, MDR_RAM13, MDR_RAM12, MDR_RAM11, MDR_RAM10, MDR_RAM9, MDR_RAM8, 
	MDR_RAM7,  MDR_RAM6,  MDR_RAM5,  MDR_RAM4,  MDR_RAM3,  MDR_RAM2,  MDR_RAM1, MDR_RAM0, 
	// from memory
	MEMMDR15, MEMMDR14, MEMMDR13, MEMMDR12, MEMMDR11, MEMMDR10, MEMMDR9, MEMMDR8,
	MEMMDR7,  MEMMDR6,  MEMMDR5,  MEMMDR4,  MEMMDR3,  MEMMDR2,  MEMMDR1, MEMMDR0,
	// from trace
	TRACEMDR15, TRACEMDR14, TRACEMDR13, TRACEMDR12, TRACEMDR11, TRACEMDR10, TRACEMDR9, TRACEMDR8,
	TRACEMDR7,  TRACEMDR6,  TRACEMDR5,  TRACEMDR4,  TRACEMDR3,  TRACEMDR2,  TRACEMDR1, TRACEMDR0,
	// from status
	STATEMDR15, STATEMDR14, STATEMDR13, STATEMDR12, STATEMDR11, STATEMDR10, STATEMDR9, STATEMDR8,
	STATEMDR7,  STATEMDR6,  STATEMDR5,  STATEMDR4,  STATEMDR3,  STATEMDR2,  STATEMDR1, STATEMDR0,
	// from break
	BRKMDR15, BRKMDR14, BRKMDR13, BRKMDR12, BRKMDR11, BRKMDR10, BRKMDR9, BRKMDR8,
	BRKMDR7,  BRKMDR6,  BRKMDR5,  BRKMDR4,  BRKMDR3,  BRKMDR2,  BRKMDR1, BRKMDR0,
	// from host if
	HOSTIFMDR15, HOSTIFMDR14, HOSTIFMDR13, HOSTIFMDR12, HOSTIFMDR11, HOSTIFMDR10, HOSTIFMDR9, HOSTIFMDR8,
	HOSTIFMDR7,  HOSTIFMDR6,  HOSTIFMDR5,  HOSTIFMDR4,  HOSTIFMDR3,  HOSTIFMDR2,  HOSTIFMDR1, HOSTIFMDR0,
	// from dflashemu
	DFMDR15, DFMDR14, DFMDR13, DFMDR12, DFMDR11, DFMDR10, DFMDR9, DFMDR8,
	DFMDR7,  DFMDR6,  DFMDR5,  DFMDR4,  DFMDR3,  DFMDR2,  DFMDR1, DFMDR0,
	// etc.
	SLDFLASH
	);

	output	MDR_RAM15, MDR_RAM14, MDR_RAM13, MDR_RAM12, MDR_RAM11, MDR_RAM10, MDR_RAM9, MDR_RAM8, 
		MDR_RAM7,  MDR_RAM6,  MDR_RAM5,  MDR_RAM4,  MDR_RAM3,  MDR_RAM2,  MDR_RAM1, MDR_RAM0;
	input	MEMMDR15, MEMMDR14, MEMMDR13, MEMMDR12, MEMMDR11, MEMMDR10, MEMMDR9, MEMMDR8,
		MEMMDR7,  MEMMDR6,  MEMMDR5,  MEMMDR4,  MEMMDR3,  MEMMDR2,  MEMMDR1, MEMMDR0;
	input	TRACEMDR15, TRACEMDR14, TRACEMDR13, TRACEMDR12, TRACEMDR11, TRACEMDR10, TRACEMDR9, TRACEMDR8,
		TRACEMDR7,  TRACEMDR6,  TRACEMDR5,  TRACEMDR4,  TRACEMDR3,  TRACEMDR2,  TRACEMDR1, TRACEMDR0;
	input	STATEMDR15, STATEMDR14, STATEMDR13, STATEMDR12, STATEMDR11, STATEMDR10, STATEMDR9, STATEMDR8,
		STATEMDR7,  STATEMDR6,  STATEMDR5,  STATEMDR4,  STATEMDR3,  STATEMDR2,  STATEMDR1, STATEMDR0;
	input	BRKMDR15, BRKMDR14, BRKMDR13, BRKMDR12, BRKMDR11, BRKMDR10, BRKMDR9, BRKMDR8,
		BRKMDR7,  BRKMDR6,  BRKMDR5,  BRKMDR4,  BRKMDR3,  BRKMDR2,  BRKMDR1, BRKMDR0;
	input	HOSTIFMDR15, HOSTIFMDR14, HOSTIFMDR13, HOSTIFMDR12, HOSTIFMDR11, HOSTIFMDR10, HOSTIFMDR9, HOSTIFMDR8,
		HOSTIFMDR7,  HOSTIFMDR6,  HOSTIFMDR5,  HOSTIFMDR4,  HOSTIFMDR3,  HOSTIFMDR2,  HOSTIFMDR1, HOSTIFMDR0;
	input	DFMDR15, DFMDR14, DFMDR13, DFMDR12, DFMDR11, DFMDR10, DFMDR9, DFMDR8,
		DFMDR7,  DFMDR6,  DFMDR5,  DFMDR4,  DFMDR3,  DFMDR2,  DFMDR1, DFMDR0;
        input   SLDFLASH;

	wire [15:0]	mdr, mdr1, mdr2, mdr3, mdr4, mdr5, mdr6;

	assign	{MDR_RAM15, MDR_RAM14, MDR_RAM13, MDR_RAM12, MDR_RAM11, MDR_RAM10, MDR_RAM9, MDR_RAM8, 
		MDR_RAM7,  MDR_RAM6,  MDR_RAM5,  MDR_RAM4,  MDR_RAM3,  MDR_RAM2,  MDR_RAM1, MDR_RAM0} = mdr;

	assign	mdr1 = {MEMMDR15, MEMMDR14, MEMMDR13, MEMMDR12, MEMMDR11, MEMMDR10, MEMMDR9, MEMMDR8,
			MEMMDR7,  MEMMDR6,  MEMMDR5,  MEMMDR4,  MEMMDR3,  MEMMDR2,  MEMMDR1, MEMMDR0};
	assign	mdr2 = {TRACEMDR15, TRACEMDR14, TRACEMDR13, TRACEMDR12, TRACEMDR11, TRACEMDR10, TRACEMDR9, TRACEMDR8,
			TRACEMDR7,  TRACEMDR6,  TRACEMDR5,  TRACEMDR4,  TRACEMDR3,  TRACEMDR2,  TRACEMDR1, TRACEMDR0};
	assign	mdr3 = {STATEMDR15, STATEMDR14, STATEMDR13, STATEMDR12, STATEMDR11, STATEMDR10, STATEMDR9, STATEMDR8,
			STATEMDR7,  STATEMDR6,  STATEMDR5,  STATEMDR4,  STATEMDR3,  STATEMDR2,  STATEMDR1, STATEMDR0};
	assign	mdr4 = {BRKMDR15, BRKMDR14, BRKMDR13, BRKMDR12, BRKMDR11, BRKMDR10, BRKMDR9, BRKMDR8,
			BRKMDR7,  BRKMDR6,  BRKMDR5,  BRKMDR4,  BRKMDR3,  BRKMDR2,  BRKMDR1, BRKMDR0};
	assign	mdr5 = {HOSTIFMDR15, HOSTIFMDR14, HOSTIFMDR13, HOSTIFMDR12, HOSTIFMDR11, HOSTIFMDR10, HOSTIFMDR9, HOSTIFMDR8,
			HOSTIFMDR7,  HOSTIFMDR6,  HOSTIFMDR5,  HOSTIFMDR4,  HOSTIFMDR3,  HOSTIFMDR2,  HOSTIFMDR1, HOSTIFMDR0};
	assign	mdr6 = {DFMDR15, DFMDR14, DFMDR13, DFMDR12, DFMDR11, DFMDR10, DFMDR9, DFMDR8,
			DFMDR7,  DFMDR6,  DFMDR5,  DFMDR4,  DFMDR3,  DFMDR2,  DFMDR1, DFMDR0};

	assign mdr = {~SLDFLASH & mdr1[15] , ~SLDFLASH & mdr1[14] , ~SLDFLASH & mdr1[13] , ~SLDFLASH & mdr1[12] , // When DataFlash read, IRAM should not out.
		      ~SLDFLASH & mdr1[11] , ~SLDFLASH & mdr1[10] , ~SLDFLASH & mdr1[9]  , ~SLDFLASH & mdr1[8]  ,
		      ~SLDFLASH & mdr1[7]  , ~SLDFLASH & mdr1[6]  , ~SLDFLASH & mdr1[5]  , ~SLDFLASH & mdr1[4]  , 
		      ~SLDFLASH & mdr1[3]  , ~SLDFLASH & mdr1[2]  , ~SLDFLASH & mdr1[1]  , ~SLDFLASH & mdr1[0]  }
	             | mdr2 | mdr3 | mdr4 | mdr5 | mdr6;

endmodule


module add_1695(DIN,DIN2,DIN3,DIN4,DIN5,DIN6,DOUT,DOUT4);
   input DIN;
   input [2:0]  DIN2;
   input [2:0]	DIN3;
   input 		DIN5;
   input [2:0] 	DIN6;
	
   
   output DOUT;
   input [2:0] DIN4;
   output DOUT4;   
endmodule // add_1695

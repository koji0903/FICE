module ConnectB(I);
   input I;   
endmodule // ConnectA

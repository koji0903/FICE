module port8_ICE(SPAD,PTTL,PTTL2,rst_b,SCANCLK)/*synthesis syn_black_box*/;
   inout SPAD;   
   input PTTL;
   input PTTL2;
   input SCANCLK;
   
   output rst_b;

endmodule // port8

module SubMod_Replace(a,add_in_port,c,d);
   input a;
   
//   input [3:0] b;
   input 	   add_in_port;
   
   output c;
   output d;   
endmodule